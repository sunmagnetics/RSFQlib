* Author: L. Schindler
* Version: 1.1.40
* Last modification date: 30 January 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

* Ports 			IN CLK OUT	
.subckt LSmitll_DFFT a clk q
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01rx1=0.7938
.param B01rx2=0.9061
.param B01tx1=3.0271
.param B02rx2=0.9638
.param B1=1.4278
.param B2=1.4988 
.param B3=0.9602 
.param B4=1.6952 
.param B5=1.1735 
.param B6=1.3640 
.param B7=1.5000 
.param IB01rx1=0.000115456 
.param IB01rx2=0.000101889 
.param IB01tx1=0.000181403 
.param IB1=0.0001204024 
.param IB2=6.34786e-005 
.param IB3=0.000153633 
.param IB4=0.00016173 
.param L01rx1=1.4067e-012 
.param L01rx2=1.2310e-012 
.param L02rx1=3.2947e-012 
.param L02rx2=2.4404e-012 
.param L02tx1=1.8040e-012 
.param L03rx2=3.6494e-012 
.param L1=1.1285e-012 
.param L2a=5.4028e-013 
.param L2b=1.6029e-012 
.param L3=9.4537e-013 
.param L3a=1.1141e-012 
.param L4=4.4401e-012 
.param L5a=3.6349e-012 
.param L5b=5.9394e-013 
.param L6=1.3233e-012 
.param L7=1.9079e-012 
.param L8=1.7976e-012 
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01rx2=(RB01rx2/Rsheet)*Lsheet
.param LRB01tx1=(RB01tx1/Rsheet)*Lsheet
.param LRB02rx2=(RB02rx2/Rsheet)*Lsheet
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param RB01rx2=B0Rs/B01rx2
.param RB01rx1=B0Rs/B01rx1
.param RB01tx1=B0Rs/B01tx1
.param RB02rx2=B0Rs/B02rx2
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
B01rx1 10 32 54 jjmit area=B01rx1
B01rx2 4 18 49 jjmit area=B01rx2
B01tx1 15 47 59 jjmit area=B01tx1
B02rx2 5 21 50 jjmit area=B02rx2
B1 11 35 55 jjmit area=B1
B2 8 9 53 jjmit area=B2
B3 12 38 56 jjmit area=B3
B4 13 41 57 jjmit area=B4
B5 7 13 52 jjmit area=B5
B6 6 24 51 jjmit area=B6
B7 14 44 58 jjmit area=B7
IB01rx1 0 34 pwl(0 0 5p IB01rx1)
IB01rx2 0 20 pwl(0 0 5p IB01rx2)
IB01tx1 0 46 pwl(0 0 5p IB01tx1)
IB1 0 37 pwl(0 0 5p IB1)
IB2 0 40 pwl(0 0 5p IB2)
IB3 0 43 pwl(0 0 5p IB3)
IB4 0 23 pwl(0 0 5p IB4)
L01rx1 a 10 L01rx1
L01rx2 clk 4 L01rx2
L02rx1 10 27 L02rx1
L02rx2 4 16 L02rx2
L02tx1 15 31 L02tx1
L03rx2 16 5 L03rx2
L1 27 11 L1
L2a 11 28 L2a
L2b 28 8 L2b
L3 12 29 L3
L3a 9 12 L3a
L4 29 13 L4
L5a 13 30 L5a
L5b 30 14 L5b
L6 14 15 L6
L7 6 7 L7
L8 5 6 L8
LIB01tx1 15 46 0.2p
LIB2 29 40 0.2p
LIB3 30 43 0.2p
LP01rx1 32 0 0.34p
LP01rx2 18 0 0.34p
LP01tx1 47 0 5e-14
LP02rx2 21 0 0.06p
LP1 35 0 0.2p
LP3 38 0 0.2p
LP4 41 0 0.2p
LP6 24 0 0.2p
LPB7 44 0 0.2p
LPIB1 28 37 0.2p
LPIB4 6 23 0.2p
LPR01rx1 27 34 0.2p
LPR01rx2 16 20 2e-13
LRB01rx1 33 0 LRB01rx1
LRB01rx2 19 0 LRB01rx2
LRB01tx1 48 0 LRB01tx1
LRB02rx2 22 0 LRB02rx2
LRB1 36 0 LRB1
LRB2 26 9 LRB2
LRB3 39 0 LRB3
LRB4 42 0 LRB4
LRB5 25 13 LRB5
LRB6 17 0 LRB6
LRB7 45 0 LRB7
RB01rx1 10 33 RB01rx1
RB01rx2 4 19 RB01rx2
RB01tx1 15 48 RB01tx1
RB02rx2 5 22 RB02rx2
RB1 11 36 RB1
RB2 8 26 RB2
RB3 12 39 RB3
RB4 13 42 RB4
RB5 7 25 RB5
RB6 6 17 RB6
RB7 14 45 RB7
RINStx1 31 q 1.36
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.ends LSmitll_DFFT