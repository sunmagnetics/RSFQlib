* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===
* Back-annotated simulation file written by InductEx v.6.0.4 on 14-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 11 June 2021
* Last modification by: L. Schindler
* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University
* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:
* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.
* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.
*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za
*$Ports    a q
.subckt LSMITLL_BUFF a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param B2=IC
.param B3=IC
.param B4=IC
.param IB1=B1*Ic0*BiasCoef
.param IB2=B2*Ic0*0.95
.param IB3=B3*Ic0*0.95
.param IB4=B4*Ic0*BiasCoef
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)
.param L4=Phi0/(2*B3*Ic0)
.param L5=Phi0/(4*IC*Ic0)
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP4=LP
B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 7 8 jjmit area=B3
B4 10 11 jjmit area=B4
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 9 pwl(0 0 5p IB3)
IB4 0 12 pwl(0 0 5p IB4)
L1 a 1 2.057E-12
L2 1 4 4.026E-12
L3 4 7 4.155E-12
L4 7 10 4.057E-12
L5 10 q 2.057E-12
LP1 2 0 5.283E-13
LP2 5 0 5.327E-13
LP3 8 0 5.084E-13
LP4 11 0 5.269E-13
LB1 1 3 LB1
LB2 4 6 LB2
LB3 7 9 LB3
LB4 10 12 LB4
RB1 1 101 RB1
RB2 4 104 RB2
RB3 7 107 RB3
RB4 10 110 RB4
LRB1 101 0 LRB1
LRB2 104 0 LRB2
LRB3 107 0 LRB3
LRB4 110 0 LRB4
.ends
* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 11
b1   1  2  jjmitll100 area=2.25
b2   3  4  jjmitll100 area=2.25
b3   5  6  jjmitll100 area=2.5
ib1  0  2  pwl(0 0 5p 275ua)
ib2  0  5  pwl(0 0 5p 175ua)
l1   8  7  1p
l2   7  0  3.9p
l3   7  1  0.6p
l4   2  3  1.1p
l5   3  5  4.5p
l6   5  11 2p
lp2  4  0  0.2p
lp3  6  0  0.2p
lrb1 9  2  1p
lrb2 10 4  1p
lrb3 12 6  1p
rb1  1  9  4.31
rb2  3  10 4.31
rb3  5  12 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.2p
.param ic=2.5
.param lptl=2p
.param lb=2p
.param biascoef=0.7
.param b1=ic
.param b2=ic
.param ib1=(b1+b2)*ic0*biascoef
.param lb1=lb
.param l1=phi0/(4*b1*ic0)
.param l2=phi0/(4*b1*ic0)
.param l3=phi0/(4*b1*ic0)
.param l4=phi0/(4*b2*ic0)
.param rb1=2.743962
.param rb2=2.743962
.param lrb1=1.750339e-12
.param lrb2=1.750339e-12
.param lp1=lp
.param lp2=lp
b1 1 2 jjmit area=b1
b2 6 7 jjmit area=b2
ib1 0 5 pwl(0 0 5p ib1)
l1 a 1 l1
l2 1 4 l2
l3 4 6 l3
l4 6 q l4
lp1 2 0 lp1
lp2 7 0 lp2
lb1 5 4 lb1
rb1 1 3 rb1
rb2 6 8 rb2
lrb1 3 0 lrb1
lrb2 8 0 lrb2
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.2p
.param ic=2.5
.param lptl=2p
.param lb=2p
.param biascoef=0.7
.param b1=ic
.param b2=ic
.param ib1=(b1+b2)*ic0*biascoef
.param lb1=lb
.param l1=phi0/(4*b1*ic0)
.param l2=phi0/(4*b1*ic0)
.param l3=phi0/(4*b1*ic0)
.param l4=phi0/(4*b2*ic0)
.param rb1=2.743962
.param rb2=2.743962
.param lrb1=1.750339e-12
.param lrb2=1.750339e-12
.param lp1=lp
.param lp2=lp
b1 1 2 jjmit area=b1
b2 6 7 jjmit area=b2
ib1 0 5 pwl(0 0 5p ib1)
l1 a 1 l1
l2 1 4 l2
l3 4 6 l3
l4 6 q l4
lp1 2 0 lp1
lp2 7 0 lp2
lb1 5 4 lb1
rb1 1 3 rb1
rb2 6 8 rb2
lrb1 3 0 lrb1
lrb2 8 0 lrb2
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  1
r1 1 0 2
.ENDS SINKCELL
* ===== MAIN =====
I_a 0 1 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa SOURCECELL 1 2
XLOADINa LOADINCELL 2 3
XLOADOUTq LOADOUTCELL 4 5
XSINKOUTq SINKCELL 5
XDUT lsmitll_buff 3 4
.tran 0.025p 1000p 0
.print i(L1.XDUT) p(B1.XDUT) i(L5.XDUT) p(B4.XDUT)
.end
