* Author: L. Schindler
* Version: 2.1
* Last modification date: 26 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			  a q0 q1
.subckt LSMITLL_SPLITT a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param Lptl=2p
.param BiasCoef=0.7
.param RD=1.36
.param B1=ICreceive
.param B2=IC
.param B3=ICtrans
.param B4=ICtrans
.param IB1=BiasCoef*(B1+B2)*Ic0
.param IB2=BiasCoef*B3*Ic0
.param IB3=BiasCoef*B4*Ic0
.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))/2
.param L3=(Phi0/(2*B1*Ic0))/2
.param L4=(Phi0/(2*B2*Ic0))/2
.param L5=(Phi0/(2*B2*Ic0))/2
.param L6=Lptl
.param L7=(Phi0/(2*B2*Ic0))/2
.param L8=Lptl
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 8 pwl(0 0 5p IB2)
IB3 0 11 pwl(0 0 5p IB3)
B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 8 9 jjmit area=B3
B4 11 12 jjmit area=B4
L1 a 2 L1
L2 2 4 L2
L3 4 5 L3
L4 5 7 L4
L5 7 8 L5
L6 8 10 L6
L7 7 11 L7
L8 11 13 L8
LP1 3 0 0.2p
LP2 6 0 0.2p
LP3 9 0 0.2p
LP4 12 0 0.2p
RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 8 108 RB3
LRB3 108 0 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
RD1 13 q0 RD
RD2 10 q1 RD
.ends