* Back-annotated simulation file written by InductEx v.6.0.4 on 30-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 11 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports  				a  q
.subckt LSmitll_bufft  a  q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param RD=1.36
.param LB=0.2p
.param Lptl=2p
.param LP=0.5p

.param B1=2.0
.param B2=2.5
.param B3=2.5
.param IB1=168u
.param IB2=340u
.param LB1=LB
.param LB2=LB
.param L1=Lptl
.param L2=6.2p
.param L3=2.07p
.param L4=2.07p
.param L5=Lptl
.param LP1=LP
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 6 7 jjmit area=B2
B3 11 12 jjmit area=B3
IB1 0 5 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
L1 a 2 2.727E-12
L2 2 6 6.22E-12  
L3 6 9 2.06E-12
L4 9 11 2.051E-12
L5 11 14 2.041E-12
RD 14 q RD
LP1 3 0 5.275E-13
LP2 7 0 5.212E-13
LP3 12 0 5.126E-13
RB1 2 4 RB1
RB2 6 8 RB2
RB3 11 13 RB3
LRB1 4 0 LRB1
LRB2 8 0 LRB2
LRB3 13 0 LRB3
LB1 2 5 2.883E-12
LB2 9 10 2.393E-12
.ends