* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 2 June 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_Always0_async_v2p1.cir
.endc

L1 a 1 [L1]
L2 1 4 [L2]
L3 5 6 [L3]
L4 6 q [L4]

LB1 1 3 [LB1]
LB2 6 8 [LB2]
LP1 2 0 [LP1]
LP2 7 0 [LP2]

* Ports
P1 a 0
P2 q 0
J1 1 2 250
J2 6 7 250
PB1 3 0
PB2 8 0
PR1 4 0
PR2 5 0
.ends