* Adapted from Fluxonics SDQDC_v5
* Author: L. Schindler
* Version: 2.1
* Last modification date: 23 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports a q
.subckt LSmitll_SFQDC a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12
.param LB=2p
.param LP=0.5p

.param B1=3.25
.param B2=2.00
.param B3=1.50
.param B4=3.00
.param B5=1.75
.param B6=1.50
.param B7=1.50
.param B8=2.00

.param IB1=280u
.param IB2=150u
.param IB3=220u
.param IB4=80u

.param L1=1.522p
.param L3=0.827p
.param L4=1.12884p
.param L5=1.11098p
.param L5b=3.216p
.param L6=5.94p
.param L10=0.215p
.param L19=0.954p
.param L13=3.699p
.param L18=2.010p
.param L17=1.510p
.param LR1=0.91p
.param R1=0.375

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LP1=LP
.param LP4=LP
.param LP5=LP
.param LP7=LP
.param LP8=LP

B1 2 4 jjmit area=B1
B2 7 10 jjmit area=B2
B3 6 8 jjmit area=B3
B4 10 11 jjmit area=B4
B5 8 15 jjmit area=B5
B6 17 18 jjmit area=B6
B7 20 21 jjmit area=B7
B8 24 25 jjmit area=B8

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 19 pwl(0 0 5p IB3)
IB4 0 23 pwl(0 0 5p IB4)

LB1 2 3 LB1
LB2 8 9 LB2
LB3 18 19 LB3
LB4 22 23 LB4

L1 a 2 L1
L3 2 5 L3
L4 5 6 L4
L5 5 7 L5
L5B 10 12 L5B
L6 8 12 L6
L10 12 17 L10
L13 20 22 L13
L17 24 q L17
L18 22 24 L18
L19 18 20 L19

LR1 12 13 LR1
R1 13 0 R1

LP1 4 0 LP1
LP4 11 0 LP4
LP5 15 0 LP5
LP7 21 0 LP7
LP8 25 0 LP8

RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 7 107 RB2
LRB2 107 10 LRB2
RB3 6 106 RB3
LRB3 106 8 LRB3
RB4 10 110 RB4
LRB4 110 0 LRB4
RB5 8 108 RB5
LRB5 108 0 LRB5
RB6 17 117 RB6
LRB6 117 18 LRB6
RB7 20 120 RB7
LRB7 120 0 LRB7
RB8 24 124 RB8
LRB8 124 0 LRB8
.ends