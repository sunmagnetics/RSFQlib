VERSION 5.8 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.01 ;

CLEARANCEMEASURE EUCLIDEAN ;

USEMINSPACING OBS ON ;

SITE CoreSite
	CLASS CORE ;
	SIZE 1 BY 160 ;
END CoreSite

LAYER M1
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M1

LAYER via1
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via1

LAYER M2
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M2

LAYER via2
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via2

LAYER M3
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M3

LAYER via3
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via3

LAYER M4
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M4

LAYER via4
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via4

LAYER M5
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M5

LAYER OVERLAP
	TYPE OVERLAP ;
END OVERLAP

VIA VIA12 DEFAULT
	LAYER M1 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via1 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M2 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA12

VIA VIA23 DEFAULT
	LAYER M2 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via2 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M3 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA23

VIA VIA34 DEFAULT
	LAYER M3 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via3 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M4 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA34

VIA VIA45 DEFAULT
	LAYER M4 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via4 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M5 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA45

MACRO PAD
	CLASS CORE ;
	ORIGIN 0.0 0.0 ;
	SIZE 100.0 BY 120.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER M1 ;
				RECT 27.0 12.5 73.0 107.5 ;
			LAYER M5 ;
				RECT 27.0 12.5 73.0 107.5 ;
		END
	END a
END PAD

MACRO THmitll_ALWAYS0T_ASYNC
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 32.8 7.2 37.2 ;
		END
	END a
END THmitll_ALWAYS0T_ASYNC

MACRO THmitll_ALWAYS0T_ASYNC_NOA
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
END THmitll_ALWAYS0T_ASYNC_NOA

MACRO THmitll_ALWAYS0T_SYNC
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 32.8 7.2 37.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 52.8 7.2 57.2 ;
		END
	END a
END THmitll_ALWAYS0T_SYNC

MACRO THmitll_ALWAYS0T_SYNC_NOA
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 32.8 7.2 37.2 ;
		END
	END clk
END THmitll_ALWAYS0T_SYNC_NOA

MACRO THmitll_AND2T
	CLASS CORE ;
	SIZE 50.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 62.8 17.2 67.2 ;
		END
	END a
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END clk
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 42.8 22.8 47.2 27.2 ;
		END
	END q
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 42.8 12.8 47.2 17.2 ;
		END
	END b
END THmitll_AND2T

MACRO THmitll_BUFFT
	CLASS CORE ;
	SIZE 20.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 2.8 17.2 7.2 ;
		END
	END q
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 42.8 17.2 47.2 ;
		END
	END a
END THmitll_BUFFT

MACRO THmitll_DCSFQ-PTLTX
	CLASS CORE ;
	SIZE 20.05 BY 70.0 ;
	ORIGIN -0.05 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
END THmitll_DCSFQ-PTLTX

MACRO THmitll_DFFT
	CLASS CORE ;
	SIZE 30.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END a
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 22.8 2.8 27.2 7.2 ;
		END
	END clk
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 22.8 62.8 27.2 67.2 ;
		END
	END q
END THmitll_DFFT

MACRO THmitll_JTLT
	CLASS CORE ;
	SIZE 20.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 2.8 17.2 7.2 ;
		END
	END q
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 32.8 17.2 37.2 ;
		END
	END a
END THmitll_JTLT

MACRO THmitll_MERGET
	CLASS CORE ;
	SIZE 50.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 42.8 32.8 47.2 37.2 ;
		END
	END q
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 42.8 62.8 47.2 67.2 ;
		END
	END b
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 2.8 17.2 7.2 ;
		END
	END a
END THmitll_MERGET

MACRO THmitll_NDROT
	CLASS CORE ;
	SIZE 50.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 42.8 62.8 47.2 67.2 ;
		END
	END b
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END a
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 22.8 7.2 27.2 ;
		END
	END clk
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 2.8 37.2 7.2 ;
		END
	END q
END THmitll_NDROT

MACRO THmitll_NOTT
	CLASS CORE ;
	SIZE 40.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END a
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 32.8 62.8 37.2 67.2 ;
		END
	END clk
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 2.8 37.2 7.2 ;
		END
	END q
END THmitll_NOTT

MACRO THmitll_OR2T
	CLASS CORE ;
	SIZE 40.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END b
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 2.8 37.2 7.2 ;
		END
	END q
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 32.8 62.8 37.2 67.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END a
END THmitll_OR2T

MACRO THmitll_SPLITT
	CLASS CORE ;
	SIZE 30.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q1
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 22.8 12.8 27.2 17.2 ;
		END
	END q1
	PIN q0
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 22.8 22.8 27.2 27.2 ;
		END
	END q0
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END a
END THmitll_SPLITT

MACRO THmitll_XORT
	CLASS CORE ;
	SIZE 50.0 BY 70.0 ;
	ORIGIN -0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END a
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 42.8 62.8 47.2 67.2 ;
		END
	END b
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 2.8 37.2 7.2 ;
		END
	END q
END THmitll_XORT

END LIBRARY
