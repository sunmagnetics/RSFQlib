* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

*$Ports 			  a b q
.subckt LSmitll_MERGET a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01rx1=0.88429 
.param B01tx1=0.842106 
.param B1=1.45438 
.param B2=0.960422 
.param B5=0.805138 
.param IB01rx1=0.000106334 
.param IB01tx1=5.04979e-5 
.param IB1=0.000186124 
.param L01rx1=2e-012 
.param L02rx1=1.27924e-012 
.param L02tx1=4.81637e-012 
.param L1=1.75737e-012 
.param L2=2e-012 
.param L6=2.22418e-012 
.param L7=8.49377e-012 
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01rx2=(RB01rx2/Rsheet)*Lsheet
.param LRB01tx1=(RB01tx1/Rsheet)*Lsheet
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param RB01rx1=B0Rs/B01rx1
.param RB01rx2=B0Rs/B01rx1
.param RB01tx1=B0Rs/B01tx1
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B1
.param RB4=B0Rs/B2
.param RB5=B0Rs/B5
B01rx1 6 18  jjmit area=B01rx1
B01rx2 13 32  jjmit area=B01rx1
B01tx1 10 28  jjmit area=B01tx1
B1 7 20  jjmit area=B1
B2 4 5  jjmit area=B2
B3 14 34  jjmit area=B1
B4 11 12  jjmit area=B2
B5 9 26  jjmit area=B5
IB01rx1 0 15 pwl(0 0 5p IB01rx1)
IB01rx2 0 24 pwl(0 0 5p IB01rx1)
IB01tx1 0 23 pwl(0 0 5p IB01tx1)
IB1 0 22 pwl(0 0 5p IB1)
L01rx1 a 6 L01rx1
L01rx2 b 13 L01rx1
L02rx1 6 16 L02rx1
L02rx2 13 30 L02rx1
L02tx1 10 25 L02tx1
L1 16 7 L1
L2 5 8 L2
L3 30 14 L1
L12 23 10 0.2p
L16 24 30 0.2p
L1b 7 4 1p
L25 28 0 0.05p
L29 34 0 0.2p
L3b 14 11 1p
L4 12 8 L2
L6 8 9 L6
L7 9 10 L7
LP01rx1 18 0 0.34p
LP01rx2 32 0 0.34p
LP1 20 0 0.2p
LP5 26 0 0.2p
LPR01rx1 15 16 0.2p
LPR1 22 8 0.2p
LRB01rx1 19 0 LRB01rx1
LRB01rx2 33 0 LRB01rx2
LRB01tx1 29 0 LRB01tx1
LRB1 21 0 LRB1
LRB2 17 5 LRB2
LRB3 35 0 LRB3
LRB4 31 12 LRB4
LRB5 27 0 LRB5
R3 25 q 1.36
RB01rx2 13 33 RB01rx2
RB01rx1 6 19 RB01rx1
RB01tx1 10 29 RB01tx1
RB1 7 21 RB1
RB2 4 17 RB2
RB3 14 35 RB3
RB4 11 31 RB4
RB5 9 27 RB5
.ends