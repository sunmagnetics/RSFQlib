* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 23 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_ALWAYS0_ASYNC_v3p0_base.cir
.endc

L1 a 1 2.0678p [L1]
L2 1 4 4.1357p [L2]
L3 5 6 4.1357p [L3]
L4 6 q 2.0678p [L4]

LB1 1 3 [LB1]
LB2 6 8 [LB2]

LP1 2 0 [LP1]
LP2 7 0 [LP2]

* Ports
P1 a 0
P2 q 0

J1 1 2 250u
J2 6 7 250u

PB1 3 0
PB2 8 0

PR1 4 0
PR2 5 0

.ends