* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/11.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 10 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	b	q
.subckt THmitll_MERGET a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=1.6
.param B2=1.10
.param B3=2.61
.param B4=1.56
.param B5=1.6
.param B6=1.10
.param B7=2.61
.param B8=1.56
.param B9=2.5

.param IB1=112u
.param IB2=170u
.param IB3=112u
.param IB4=170u
.param IB5=171u
.param IB6=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB

.param L1=Lptl
.param L2=8.8600p
.param L3=2.4587p
.param L4=1.5077p
.param L5=Lptl
.param L6=8.8600p
.param L7=2.4587p
.param L8=1.5077p
.param L9=1.0056p
.param L10=Lptl

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP9=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 7 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 14 15 jjmit  area=B6 
B7 17 18 jjmit  area=B7 
B8 17 19 jjmit  area=B8 
B9 21 22 jjmit  area=B9 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 16 pwl(0 0 5p IB4)
IB5 0 20 pwl(0 0 5p IB5)
IB6 0 23 pwl(0 0 5p IB6)

LB1 3 1 2.504E-012 
LB2 6 4 7.477E-013 
LB3 13 11 3.72E-012 
LB4 16 14 2.115E-012 
LB5 20 10 1.701E-012 
LB6 23 21 1.272E-012 

L1 a 1 1.299E-012 
L2 1 4 8.804E-012 
L3 4 7 2.465E-012 
L4 9 10 1.51E-012 
L5 b 11 1.373E-012 
L6 11 14 8.866E-012 
L7 14 17 2.459E-012 
L8 19 10 1.516E-012 
L9 10 21 1.002E-012 
L10 21 24 7.408E-013
 
RD 24 q RD  

LP1 2 0 4.76E-013 
LP2 5 0 4.103E-013 
LP3 8 0 4.056E-013 
LP5 12 0 3.991E-013 
LP6 15 0 5.058E-013 
LP7 18 0 4.187E-013 
LP9 22 0 3.717E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 7 109 RB4  
LRB4 109 9 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 14 114 RB6  
LRB6 114 0 LRB6 
RB7 17 117 RB7  
LRB7 117 0 LRB7 
RB8 17 119 RB8  
LRB8 119 19 LRB8 
RB9 21 121 RB9  
LRB9 121 0 LRB9 

.ends
