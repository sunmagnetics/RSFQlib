* Author: L. Schindler
* Version: 2.1
* Last modification date: 29 March 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_OR2_v2p1_base.cir
.endc

* Inductors
L1 a 1 2.068e-12 [L1]
L2 1 4 3.23e-12 [L2]
L3 4 6 1.2E-12 [L3]
L4 b 8 2.068e-12 [L4]
L5 8 11 3.23e-12 [L5]
L6 11 13 1.2E-12 [L6]
L7 7 15 3.28e-12 [L7]
L8 16 19 7.94e-12 [L8]
L9 clk 20 2.068e-12 [L9]
L10 20 23 3.41e-12 [L10]
L11 19 25 3.53e-12 [L11]
L12 25 q 2.068e-12 [L12]

LB1 1 3 
LB2 8 10 
LB3 7 14 
LB4 16 18 
LB5 20 22 
LB6 25 27 

LP1 2 0 [LP1]
LP2 5 0 [LP2]
LP4 9 0 [LP4]
LP5 12 0 [LP5]
LP8 17 0 [LP8]
LP9 21 0 [LP9]
LP11 24 0 [LP11]
LP12 26 0 [LP12]

* Ports
P1 a 0
P2 b 0
P3 clk 0
P4 q 0

J1 1 2 250u
J2 4 5 222u
J3 6 7 186u
J4 8 9 250u
J5 11 12 222u
J6 13 7 186u
J7 15 16 228u
J8 16 17 209u
J9 20 21 250u
J10 23 19 152u
J11 19 24 160u
J12 25 26 250u

PB1 3 0
PB2 10 0
PB3 14 0
PB4 18 0
PB5 22 0
PB6 27 0
.ends