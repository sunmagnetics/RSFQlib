* Author: L. Schindler
* Version: 2.1
* Last modification date: 4 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports a b clk q
.subckt LSmitll_XOR	a	b	clk 	q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.70
.param B1=IC
.param B2=IC
.param B3=IC
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=IC/1.25
.param B8=IC
.param B9=IC/1.25
.param B10=IC
.param B11=IC
.param IB1=BiasCoef*Ic0*B1
.param IB2=BiasCoef*Ic0*B2
.param IB3=IB1
.param IB4=IB2
.param IB5=BiasCoef*Ic0*B8
.param IB6=BiasCoef*Ic0*B11
.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=1.2p
.param L4=Phi0/(B2*Ic0)
.param L5=L1
.param L6=L2
.param L7=L3
.param L8=L4
.param L9=1.2p
.param L10=Phi0/(4*IC*Ic0)
.param L11=Phi0/(2*B8*Ic0)
.param L12=Phi0/(2*B10*Ic0)
.param L13=Phi0/(4*IC*Ic0)
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 25 6 jjmit area=B3
B4 9 10 jjmit area=B4
B5 12 13 jjmit area=B5
B6 26 14 jjmit area=B6
B7 27 16 jjmit area=B7
B8 17 18 jjmit area=B8
B9 20 16 jjmit area=B9
B10 16 21 jjmit area=B10
B11 22 23 jjmit area=B11
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 11 pwl(0 0 5p IB3)
IB4 0 15 pwl(0 0 5p IB4)
IB5 0 19 pwl(0 0 5p IB5)
IB6 0 24 pwl(0 0 5p IB6)
LB1 3 1 LB
LB2 7 6 LB
LB3 11 9 LB
LB4 15 14 LB
LB5 19 17 LB
LB6 24 22 LB
L1 a 1 L1
L2 1 4 L2
L3 4 25 L3
L4 6 8 L4
L5 b 9 L5
L6 9 12 L6
L7 12 26 L7
L8 14 8 L8
L9 8 27 L9
L10 clk 17 L10
L11 17 20 L11
L12 16 22 L12
L13 22 q L13
LP1 2 0 LP
LP2 5 0 LP
LP4 10 0 LP
LP5 13 0 LP
LP8 18 0 LP
LP10 21 0 LP
LP11 23 0 LP
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 0 LRB2
RB3 4 106 RB3
LRB3 106 6 LRB3
RB4 9 109 RB4
LRB4 109 0 LRB4
RB5 12 112 RB5
LRB5 112 0 LRB5
RB6 12 114 RB6
LRB6 114 14 LRB6
RB7 8 108 RB7
LRB7 108 16 LRB7
RB8 17 117 RB8
LRB8 117 0 LRB8
RB9 20 120 RB9
LRB9 120 16 LRB9
RB10 16 116 RB10
LRB10 116 0 LRB10
RB11 22 122 RB11
LRB11 122 0 LRB11
.ends