* Author: L. Schindler
* Version: 1.1.40
* Last modification date: 09 April 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

* Ports 			IN CLK OUT	
.subckt LSmitll_NOTT a clk q
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01=1.3488 
.param B01rx1=1.2613 
.param B01rx2=1.2476 
.param B01tx1=2.8510 
.param B02=0.7718 
.param B03=1.2227 
.param B05=1.2221 
.param B06=1.0432 
.param B07=2.2139 
.param B09=1.4100 
.param B10=1.7227 
.param B11=1.4193 
.param IB01rx1=0.000146094 
.param IB01rx2=0.000181215 
.param IB01tx1=0.000187178 
.param IB02=9.6978e-05 
.param IB03=9.5221e-05 
.param IB04=0.000101564 
.param IB06=0.000108369 
.param L01=2.2847e-12
.param L01rx1=1.8571e-12 
.param L01rx2=2.1457e-12 
.param L01tx1=4.5195e-12 
.param L02rx1=4.4718e-12 
.param L02rx2=2.5468e-12 
.param L02tx1=3.4724e-12 
.param L03=6.5962e-12 
.param L04=4.2413e-13 
.param L06=3.2860e-12 
.param L07=4.9986e-13 
.param L08=8.6946e-13 
.param L09=2.8417e-13 
.param L10=7.3651e-12 
.param L12=2.6532e-12
.param L13=2.1566e-12 
.param L16=2.6117e-12 
.param L17=9.9180e-13 
.param L18=2.5842e-13 
.param L19=3.1681e-12 
.param L20=1.1676e-12 
.param L21=7.4611e-13 
.param LRB01=(RB01/Rsheet)*Lsheet
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01rx2=(RB01rx2/Rsheet)*Lsheet
.param LRB01tx1=(RB01tx1/Rsheet)*Lsheet
.param LRB02=(RB02/Rsheet)*Lsheet
.param LRB03=(RB03/Rsheet)*Lsheet
.param LRB05=(RB05/Rsheet)*Lsheet
.param LRB06=(RB06/Rsheet)*Lsheet
.param LRB07=(RB07/Rsheet)*Lsheet
.param LRB09=(RB09/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param RB01=B0Rs/B01
.param RB01rx1=B0Rs/B01rx1
.param RB01rx2=B0Rs/B01rx2
.param RB01tx1=B0Rs/B01tx1
.param RB02=B0Rs/B02
.param RB03=B0Rs/B03
.param RB05=B0Rs/B05
.param RB06=B0Rs/B06
.param RB07=B0Rs/B07
.param RB09=B0Rs/B09
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
B01 4 5 58 jjmit area=B01
B01rx1 17 49 64 jjmit area=B01rx1
B01rx2 12 37 60 jjmit area=B01rx2
B01tx1 8 29 57 jjmit area=B01tx1
B02 14 9 59 jjmit area=B02
B03 14 15 63 jjmit area=B03
B05 10 41 62 jjmit area=B05
B06 6 25 55 jjmit area=B06
B07 13 39 61 jjmit area=B07
B09 7 27 56 jjmit area=B09
B10 19 53 66 jjmit area=B10
B11 18 51 65 jjmit area=B11
IB01rx1 0 44 pwl(0 0 5p IB01rx1)
IB01rx2 0 31 pwl(0 0 5p IB01rx2)
IB01tx1 0 21 pwl(0 0 5p IB01tx1)
IB02 0 33 pwl(0 0 5p IB02)
IB03 0 32 pwl(0 0 5p IB03)
IB04 0 45 pwl(0 0 5p IB04)
IB06 0 20 pwl(0 0 5p IB06)
L01 10 4 L01
L01rx1 a 17 L01rx1
L01rx2 clk 12 L01rx2
L01tx1 7 8 L01tx1
L02rx1 17 46 L02rx1
L02rx2 12 34 L02rx2
L02tx1 8 24 L02tx1
L03 10 36 L03
L04 36 14 L04
L06 35 10 L06
L07 5 9 L07
L08 15 16 L08
L09 5 6 L09
L10 6 22 L10
L12 47 16 L12
L13 34 13 L13
L16 46 18 L16
L17 13 35 L17
L18 16 19 L18
L19 19 48 L19
L20 18 47 L20
L21 22 7 L21
LP01rx1 49 0 0.34p
LP01rx2 37 0 0.34p
LP01tx1 29 0 0.05p
LP05 41 0 0.567p
LP06 25 0 0.27p
LP07 39 0 0.328p
LP09 27 0 0.12p
LP10 53 0 0.239p
LP11 51 0 0.109p
LPR01rx1 46 44 0.2p
LPR01rx2 31 34 0.2p
LPR01tx1 21 8 0.2p
LPR02 33 36 0.023p
LPR03 32 35 0.208p
LPR04 47 45 0.216p
LPR06 20 22 0.13p
LRB01 23 5 LRB01
LRB01rx1 50 0 LRB01rx1
LRB01rx2 38 0 LRB01rx2
LRB01tx1 30 0 LRB01tx1
LRB02 9 11 LRB02
LRB03 43 15 LRB03
LRB05 42 0 LRB05
LRB06 26 0 LRB06
LRB07 40 0 LRB07
LRB09 28 0 LRB09
LRB10 54 0 LRB10
LRB11 52 0 LRB11
RB01 4 23 RB01
RB01rx1 17 50 RB01rx1
RB01rx2 12 38 RB01rx2
RB01tx1 8 30 RB01tx1
RB02 11 14 RB02
RB03 14 43 RB03
RB05 10 42 RB05
RB06 6 26 RB06
RB07 13 40 RB07
RB09 7 28 RB09
RB10 19 54 RB10
RB11 18 52 RB11
RD 48 0 3.54
RINStx1 24 q 1.36
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.ends LSmitll_NOTT