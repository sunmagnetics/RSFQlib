* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 29 July 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_BUFF_v3p0_base.cir
.endc

* Inductors
L1 a 1 2.0678p [L1]
L2 1 4 4.1357p [L2]
L3 4 7 4.1357p [L3]
L4 7 10 4.1357p [L4]
L5 10 q 2.0678p [L5]

LB1 1 3 
LB2 4 6 
LB3 7 9 
LB4 10 12 

LP1 2 0 [LP1]
LP2 5 0 [LP2]
LP3 8 0 [LP3]
LP4 11 0 [LP4]

* Ports
P1 a 0 
P2 q 0

J1 1 2 250u
J2 4 5 250u
J3 7 8 250u
J4 10 11 250u

PB1 3 0
PB2 6 0
PB3 9 0
PB4 12 0
.end