VERSION 5.8 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.01 ;

CLEARANCEMEASURE EUCLIDEAN ;

USEMINSPACING OBS ON ;

SITE CoreSite
	CLASS CORE ;
	SIZE 1 BY 160 ;
END CoreSite

LAYER M1
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M1

LAYER via1
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via1

LAYER M2
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M2

LAYER via2
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via2

LAYER M3
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M3

LAYER via3
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via3

LAYER M4
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M4

LAYER via4
	TYPE CUT ;
	SPACING 5.6 ;
	WIDTH 4.4 ;
END via4

LAYER M5
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 4.4 ;
	SPACING 5.6 ;
	SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
	SPACINGTABLE
		PARALLELRUNLENGTH 0.0
		WIDTH 0.0 0.06
		WIDTH 0.1 0.1
		WIDTH 0.75 0.25
		WIDTH 1.5 0.45 ;
	PITCH 10.0 10.0 ;
END M5

LAYER OVERLAP
	TYPE OVERLAP ;
END OVERLAP

VIA VIA12 DEFAULT
	LAYER M1 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via1 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M2 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA12

VIA VIA23 DEFAULT
	LAYER M2 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via2 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M3 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA23

VIA VIA34 DEFAULT
	LAYER M3 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via3 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M4 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA34

VIA VIA45 DEFAULT
	LAYER M4 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER via4 ;
		RECT -2.2 -2.2 2.2 2.2 ;
	LAYER M5 ;
		RECT -2.2 -2.2 2.2 2.2 ;
END VIA45

MACRO PAD
	CLASS CORE ;
	ORIGIN 0.0 0.0 ;
	SIZE 100.0 BY 120.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INOUT ;
	USE SIGNAL ;
		PORT
			LAYER M1 ;
				RECT 27.0 12.5 73.0 107.5 ;
			LAYER M5 ;
				RECT 27.0 12.5 73.0 107.5 ;
		END
	END a
END PAD

MACRO LSmitll_OR2T
	CLASS CORE ;
	SIZE 100.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 82.8 52.8 87.2 57.2 ;
		END
	END clk
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END b
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 82.8 12.8 87.2 17.2 ;
		END
	END q
END LSmitll_OR2T

MACRO LSmitll_JTLT
	CLASS CORE ;
	SIZE 40.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 52.8 7.2 57.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 12.8 37.2 17.2 ;
		END
	END q
END LSmitll_JTLT

MACRO LSmitll_PTLRX_SFQDC
	CLASS CORE ;
	SIZE 100.1 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
END LSmitll_PTLRX_SFQDC

MACRO LSmitll_MERGET
	CLASS CORE ;
	SIZE 70.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END b
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 62.8 12.8 67.2 17.2 ;
		END
	END q
END LSmitll_MERGET

MACRO LSmitll_PTLTX
	CLASS CORE ;
	SIZE 30.1 BY 70.0 ;
	ORIGIN -0.1 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 22.8 22.8 27.2 27.2 ;
		END
	END Q
END LSmitll_PTLTX

MACRO LSmitll_Always0T_sync
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 32.8 7.2 37.2 ;
		END
	END a
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END clk
END LSmitll_Always0T_sync

MACRO LSmitll_SPLITT
	CLASS CORE ;
	SIZE 50.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
	PIN q0
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 2.8 17.2 7.2 ;
		END
	END q0
	PIN q1
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 2.8 37.2 7.2 ;
		END
	END q1
END LSmitll_SPLITT

MACRO LSmitll_NDROT
	CLASS CORE ;
	SIZE 120.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN in_clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 102.8 52.8 107.2 57.2 ;
		END
	END in_clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END b
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 102.8 12.8 107.2 17.2 ;
		END
	END q
END LSmitll_NDROT

MACRO LSmitll_DFFT
	CLASS CORE ;
	SIZE 80.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 62.8 12.8 67.2 17.2 ;
		END
	END q
END LSmitll_DFFT

MACRO LSmitll_Always0T_sync
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 2.8 62.8 7.2 67.2 ;
		END
	END clk
END LSmitll_Always0T_sync

MACRO LSmitll_PTLRX
	CLASS CORE ;
	SIZE 40.1 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
END LSmitll_PTLRX

MACRO LSmitll_Always0T_async
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 32.8 7.2 37.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
END LSmitll_Always0T_async

MACRO LSmitll_Always0T_async_noA
	CLASS CORE ;
	SIZE 10.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 2.8 7.2 7.2 ;
		END
	END q
END LSmitll_Always0T_async_noA

MACRO LSmitll_AND2T
	CLASS CORE ;
	SIZE 100.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 82.8 52.8 87.2 57.2 ;
		END
	END b
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 82.8 12.8 87.2 17.2 ;
		END
	END q
END LSmitll_AND2T

MACRO LSmitll_XORT
	CLASS CORE ;
	SIZE 100.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 82.8 52.8 87.2 57.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END b
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 82.8 12.8 87.2 17.2 ;
		END
	END q
END LSmitll_XORT

MACRO LSmitll_XNORT
	CLASS CORE ;
	SIZE 90.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 72.8 12.8 77.2 17.2 ;
		END
	END Q
	PIN b
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END b
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END a
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 62.8 52.8 67.2 57.2 ;
		END
	END clk
END LSmitll_XNORT

MACRO LSmitll_NOTT
	CLASS CORE ;
	SIZE 100.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN clk
	DIRECTION INPUT ;
	USE CLOCK ;
		PORT
			LAYER M3 ;
				RECT 12.8 52.8 17.2 57.2 ;
		END
	END clk
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 12.8 12.8 17.2 17.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 82.8 12.8 87.2 17.2 ;
		END
	END q
END LSmitll_NOTT

MACRO LSmitll_BUFFT
	CLASS CORE ;
	SIZE 40.0 BY 70.0 ;
	ORIGIN 0.0 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN a
	DIRECTION INPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 2.8 52.8 7.2 57.2 ;
		END
	END a
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 32.8 12.8 37.2 17.2 ;
		END
	END q
END LSmitll_BUFFT

MACRO LSmitll_DCSFQ-PTLTX
	CLASS CORE ;
	SIZE 60.1 BY 50.0 ;
	ORIGIN -0.1 0.0 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN q
	DIRECTION OUTPUT ;
	USE SIGNAL ;
		PORT
			LAYER M3 ;
				RECT 52.8 12.8 57.2 17.2 ;
		END
	END q
END LSmitll_DCSFQ-PTLTX

END LIBRARY
