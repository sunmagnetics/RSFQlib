* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 2 June 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_Always0_sync_v2p1.cir
.endc

L1 a 1 [L1]
L2 1 4 [L2]
L3 clk 5 [L3]
L4 5 8 [L4]
L5 9 10 [L5]
L6 10 q [L6]

LB1 1 3 [LB1]
LB2 5 7 [LB2]
LB3 10 12 [LB3]
LP1 2 0 [LP1]
LP2 6 0 [LP2]
LP3 11 0 [LP3]

* Ports
P1 a 0
P2 clk 0
P3 q 0
J1 1 2 250
J2 5 6 250
J3 10 11 250
PB1 3 0
PB2 7 0
PB3 12 0
PR1 4 0
PR2 8 0
PR3 9 0
.end