* Author: L. Schindler
* Version: 2.1
* Last modification date: 27 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$ports				   a b q
.subckt LSmitll_MERGET a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.70
.param RD=1.36

.param B1=ICreceive
.param B2=IC/1.25
.param B3=IC/1.4
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=IC/1.4
.param B8=ICtrans
.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)*(B7/(B2+B7))
.param L4=L1
.param L5=L2
.param L6=L3
.param L7=Phi0/(2*B2*Ic0)*(B2/(B2+B7))
.param L8=(Phi0/(2*B7*Ic0))*(B8/(B7+B8))
.param L9=(Phi0/(2*B7*Ic0))*(B7/(B7+B8))
.param L10=Lptl
.param IB1=BiasCoef*B1*Ic0
.param IB2=IB1
.param IB3=IC*Ic0
.param IB4=BiasCoef*Ic0*(B7+B8)
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet

L1 a 1 L1
L2 1 4 L2
L3 4 6 L3
L4 b 8 L4
L5 8 11 L5
L6 11 13 L6
L7 7 15 L7
L8 15 19 L8
L9 17 19 L9
L10 19 21 L10
RD 21 q RD
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 6 7 jjmit area=B3
B4 8 9 jjmit area=B4
B5 11 12 jjmit area=B5
B6 13 7 jjmit area=B6
B7 15 16 jjmit area=B7
B8 19 20 jjmit area=B8
LP1 2 0 LP
LP2 5 0 LP
LP4 9 0 LP
LP5 12 0 LP
LP7 16 9 LP
LP8 20 0 LP
RB1 1 101 RB1
RB2 4 104 RB2
RB3 6 106 RB3
RB4 8 108 RB4
RB5 11 111 RB5
RB6 13 113 RB6
RB7 15 115 RB7
RB8 19 119 RB8
LRB1 101 0 LRB1
LRB2 104 0 LRB2
LRB3 106 7 LRB3
LRB4 108 0 LRB4
LRB5 111 0 LRB5
LRB6 113 7 LRB6
LRB7 115 0 LRB7
LRB8 119 0 LRB8
LB1 1 3 LB
LB2 8 10 LB
LB3 7 14 LB
LB4 17 18 LB
.ends