* Author: T. Hall
* Version: 3.0
* Last modification date: 24 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	clk	q
.subckt THmitll_NOTT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=ICreceive
.param B2=IC
.param B3=IC/3
.param B4=IC/3
.param B5=IC/1.4
.param B6=ICreceive
.param B7=IC
.param B8=IC/3
.param B9=IC/3
.param B10=IC

.param IB1=BiasCoef*Ic0*(B1+B2)
.param IB2=BiasCoef*Ic0*(B4+B8)
.param IB3=BiasCoef*Ic0*(B6+B7)
.param IB4=BiasCoef*B10*Ic0

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB

.param L1=Lptl
.param L2=(Phi0/(2*Ic0*B1))*(B1/(B1+B2))
.param L3=(Phi0/(2*Ic0*B1))*(B2/(B1+B2))
.param L4=Phi0/(2*B1*Ic0)
.param L5=2p
.param L6=8p
.param L7=Lptl
.param L8=(Phi0/(2*Ic0*B6))*(B6/(B6+B7))
.param L9=(Phi0/(2*Ic0*B6))*(B7/(B6+B7))
.param L10=Phi0/(2*B7*Ic0)
.param L11=2p
.param L12=8p
.param L13=Lptl

.param LP1=LP
.param LP2=LP
.param LP6=LP
.param LP7=LP
.param LP9=LP
.param LP10=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 10 11 jjmit  area=B4 
B5 12 13 jjmit  area=B5 
B6 14 15 jjmit  area=B6 
B7 18 19 jjmit  area=B7 
B8 13 20 jjmit  area=B8 
B9 11 21 jjmit  area=B9 
B10 22 23 jjmit  area=B10 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 17 pwl(0 0 5p IB3)
IB4 0 24 pwl(0 0 5p IB4)

LB1 4 3 LB1 
LB2 9 8 LB2 
LB3 17 16 LB3 
LB4 24 22 LB4 

L1 a 1 L1 
L2 1 3 L2 
L3 3 5 L3 
L4 5 7 L4 
L5 8 10 L5 
L6 8 12 L6 
L7 clk 14 L7 
L8 14 16 L8 
L9 16 18 L9 
L10 18 13 L10 
L11 11 20 L11 
L12 11 22 L12 
L13 22 25 L13 

RD 25 q RD

LP1 2 0 LP1 
LP2 6 0 LP2 
LP6 15 0 LP6 
LP7 19 0 LP7 
LP9 21 0 LP9 
LP10 23 0 LP10 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 8 LRB3 
RB4 10 110 RB4  
LRB4 110 11 LRB4 
RB5 12 112 RB5  
LRB5 112 13 LRB5 
RB6 14 114 RB6  
LRB6 114 0 LRB6 
RB7 18 118 RB7  
LRB7 118 0 LRB7 
RB8 13 113 RB8  
LRB8 113 20 LRB8 
RB9 11 111 RB9  
LRB9 111 0 LRB9 
RB10 22 122 RB10  
LRB10 122 0 LRB10 

.ends
