* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 23 June 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_Always0T_sync_v2p1_base.cir
.endc

L1 a 1 [L1]
L2 clk 2 [L2]
L3 3 q [L3]


* Ports
P1 a 0
P2 clk 0
P3 q 0
PR1 1 0
PR2 2 0
PR3 3 0
.ends