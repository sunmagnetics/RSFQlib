* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 2 June 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_DCSFQ_PTLTX_v2p1_base.cir
.endc

* Inductors
L1 1 2 [L1]
L2 2 0 3.9p [L2]
L3 2 3 0.6p [L3]
L4 4 6 1.1p [L4]
L5 6 8 4.5p [L5]
L6 8 11 4.5p [L6]
L7 11 14 3.3p [L7]
L8 14 17  [L8]
LP2 7 0 [LP2]
LP3 9 0 [LP3]
LP4 12 0 [LP4]
LP5 15 0 [LP5]
LB1 4 5 [LB1]
LB2 8 10 [LB2]
LB3 11 13 [LB3]
LB4 14 16 [LB4]
* Ports
P1 1 0
P2 17 0
PB1 5 0
PB2 10 0
PB3 13 0
PB4 16 0
J1 3 4 225u
J2 6 7 225u
J3 8 9 250u
J4 11 12 200u
J5 14 15 162u
.end