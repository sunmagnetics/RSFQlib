* Adapted from Fluxonics SDQDC_v5
* Author: L. Schindler
* Version: 3.0
* Last modification date: 13 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	q
.subckt THmitll_PTLRX-SFQDC a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=ICreceive
.param B2=IC/1.25
.param B3=3.25
.param B4=1.50
.param B5=1.75
.param B6=2.00
.param B7=3.00
.param B8=1.50
.param B9=1.50
.param B10=2.00

.param IB1=BiasCoef*Ic0*(B1+B2)
.param IB2=280u
.param IB3=150u
.param IB4=220u
.param IB5=80u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))*(B1/(B1+B2))
.param L3=(Phi0/(2*B1*Ic0))*(B2/(B1+B2))
.param L4=Phi0/(2*B2*Ic0)
.param L5=0.827p
.param L6=1.12884p
.param L7=5.94p
.param L8=1.11098p
.param L9=3.216p
.param L10=0.215p
.param L11=0.954p
.param L12=3.699p
.param L13=2.010p
.param L14=1.510p

.param LR1=0.91p
.param R1=5.74

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP5=LP
.param LP7=LP
.param LP9=LP
.param LP10=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 11 12 jjmit  area=B4 
B5 12 13 jjmit  area=B5 
B6 16 17 jjmit  area=B6 
B7 17 18 jjmit  area=B7 
B8 20 21 jjmit  area=B8 
B9 23 24 jjmit  area=B9 
B10 27 28 jjmit  area=B10 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 22 pwl(0 0 5p IB4)
IB5 0 26 pwl(0 0 5p IB5)

LB1 4 3 LB1 
LB2 9 7 LB2 
LB3 14 12 LB3 
LB4 22 21 LB4 
LB5 26 25 LB5 

L1 a 1 L1 
L2 1 3 L2 
L3 3 5 L3 
L4 5 7 L4 
L5 7 10 L5 
L6 11 10 L6 
L7 12 15 L7 
L8 10 16 L8 
L9 15 17 L9 
L10 15 20 L10 
L11 21 23 L11 
L12 23 25 L12 
L13 25 27 L13 
L14 27 q L14 

LR1 19 15 LR1 
R1 0 19 R1  

LP1 2 0 LP1 
LP2 6 0 LP2 
LP3 8 0 LP3 
LP5 13 0 LP5 
LP7 18 0 LP7 
LP9 24 0 LP9 
LP10 28 0 LP10 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 11 111 RB4  
LRB4 111 12 LRB4 
RB5 12 112 RB5  
LRB5 112 0 LRB5 
RB6 16 116 RB6  
LRB6 116 17 LRB6 
RB7 17 117 RB7  
LRB7 117 0 LRB7 
RB8 20 120 RB8  
LRB8 120 21 LRB8 
RB9 23 123 RB9  
LRB9 123 0 LRB9 
RB10 27 127 RB10  
LRB10 127 0 LRB10 

.ends
