* Circuit for InductEx extraction (excluding resistors)
* Author: T. Hall
* Version: 3.0
* Last modification date: 25 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_NOTT_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 [L1] 
L2 1 3 2.3963p [L2] 
L3 3 5 2.9984p [L3] 
L4 5 7 5.5602p [L4] 
L5 8 10 1.8403p [L5] 
L6 8 12 8.5410p [L6] 
L7 clk 14 [L7] 
L8 14 16 2.8313p [L8] 
L9 16 18 3.4874p [L9] 
L10 18 13 5.2166p [L10] 
L11 11 20 1.5349p [L11] 
L12 11 22 8.5298p [L12]
L13 22 q [L13] 

LB1 4 3 [LB1] 
LB2 9 8 [LB2] 
LB3 17 16 [LB3] 
LB4 24 22 [LB4] 

LP1 2 0 [LP1] 
LP2 6 0 [LP2] 
LP6 15 0 [LP6] 
LP7 19 0 [LP7] 
LP9 21 0 [LP9] 
LP10 23 0 [LP10] 

* Ports
P1 a 0
P2 clk 0
P3 q 0

PB1 4 0
PB2 9 0
PB3 17 0
PB4 24 0

J1 1 2 160u
J2 5 6 238u
J3 7 8 77u
J4 10 11 73u
J5 12 13 198u
J6 14 15 160u
J7 18 19 218u
J8 13 20 87u
J9 11 21 82u
J10 22 23 250u

.end