* Back-annotated simulation file written by InductEx v.6.0.4 on 2-6-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 2 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a q
.subckt LSmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1.0
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=2.25
.param B2=2.25
.param B3=2.5
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=2p
.param IB1=275u
.param IB2=175u
.param LB1=LB
.param LB2=LB
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 3 4 3.12E-12
LB2 7 9 2.281E-12
L1 a 1 1.295E-12
L2 1 0 3.904E-12
L3 1 2 5.998E-13
L4 3 5 1.095E-12
L5 5 7 4.448E-12
L6 7 q 1.334E-12
LP2 6 0 5.16E-13
LP3 8 0 4.733E-13
RB1 2 102 RB1
LRB1 102 3 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 7 107 RB3
LRB3 107 0 LRB3
.ends
