* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/08.
* Adapted from Fluxonics SDQDC_v5
* Author: L. Schindler
* Version: 3.0
* Last modification date: 4 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports 	a	q
.subckt THmitll_SFQDC a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=3.25
.param B2=1.50
.param B3=1.75
.param B4=2.00
.param B5=3.00
.param B6=1.50
.param B7=1.50
.param B8=2.00

.param IB1=280u
.param IB2=150u
.param IB3=220u
.param IB4=80u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB

.param L1=1.522p
.param L2=0.827p
.param L3=1.12884p
.param L4=5.94p
.param L5=1.11098p
.param L6=3.216p
.param L7=0.215p
.param L8=0.954p
.param L9=3.699p
.param L10=2.010p
.param L11=1.510p

.param LR1=0.91p
.param R1=0.375

.param LP1=LP
.param LP3=LP
.param LP5=LP
.param LP7=LP
.param LP8=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 6 8 jjmit  area=B3 
B4 10 11 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 14 15 jjmit  area=B6 
B7 17 18 jjmit  area=B7 
B8 21 22 jjmit  area=B8 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)

LB1 3 1 1.401E-012 
LB2 7 6 6.064E-013 
LB3 16 15 1.989E-012 
LB4 20 19 8.87E-013 

L1 a 1 1.529E-012 
L2 1 4 8.239E-013 
L3 5 4 1.124E-012 
L4 6 9 5.898E-012 
L5 4 10 1.111E-012 
L6 9 11 3.227E-012 
L7 9 14 2.138E-013 
L8 15 17 9.503E-013 
L9 17 19 3.696E-012 
L10 19 21 2.001E-012 
L11 21 q 1.496E-012 

R1 0 13 R1  
LR1 13 9 9.11E-013 

LP1 2 0 3.162E-013 
LP3 8 0 4.507E-013 
LP5 12 0 6.57E-013 
LP7 18 0 4.343E-013 
LP8 22 0 3.726E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 6 LRB2 
RB3 6 106 RB3  
LRB3 106 0 LRB3 
RB4 10 110 RB4  
LRB4 110 11 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 14 114 RB6  
LRB6 114 15 LRB6 
RB7 17 117 RB7  
LRB7 117 0 LRB7 
RB8 21 121 RB8  
LRB8 121 0 LRB8 

.ends
