* Author: L. Schindler
* Version: 3.0
* Last modification date: 30 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	b	clk	q
.subckt THmitll_XNOR a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param B3=IC/1.4
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=IC/1.4
.param B8=IC/1.25
.param B9=IC
.param B10=IC/1.4
.param B11=IC
.param B12=IC/3
.param B13=IC/3
.param B14=IC/1.4
.param B15=IC
.param B16=IC
.param B17=IC/3
.param B18=IC/3
.param B19=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=BiasCoef*Ic0*B4
.param IB3=BiasCoef*Ic0*(B3+B6)
.param IB4=BiasCoef*Ic0*B9
.param IB5=BiasCoef*Ic0*B11
.param IB6=BiasCoef*Ic0*(B14+B13)
.param IB7=BiasCoef*B15*Ic0
.param IB8=BiasCoef*B19*Ic0

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param LB8=LB

.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)
.param L4=L1
.param L5=L2
.param L6=L3
.param L7=Phi0/(2*B8*Ic0)
.param L8=Phi0/(4*IC*Ic0)
.param L9=(Phi0/(2*B9*Ic0))/2
.param L10=(Phi0/(2*B9*Ic0))/2
.param L11=Phi0/(2*B8*Ic0)
.param L12=Phi0/(2*B11*Ic0)
.param L13=2p
.param L14=4p
.param L15=(Phi0/(2*B9*Ic0))/2
.param L16=Phi0/(2*B15*Ic0)
.param L17=Phi0/(2*B16*Ic0)
.param L18=1p
.param L19=4p
.param L20=Phi0/(4*IC*Ic0)

.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP8=LP
.param LP9=LP
.param LP11=LP
.param LP15=LP
.param LP16=LP
.param LP18=LP
.param LP19=LP

.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param RB16=B0Rs/B16
.param RB17=B0Rs/B17
.param RB18=B0Rs/B18
.param RB19=B0Rs/B19

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet+LP
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet+LP
.param LRB16=(RB16/Rsheet)*Lsheet+LP
.param LRB17=(RB17/Rsheet)*Lsheet
.param LRB18=(RB18/Rsheet)*Lsheet+LP
.param LRB19=(RB19/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 4 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 11 13 jjmit  area=B6 
B7 7 15 jjmit  area=B7 
B8 16 17 jjmit  area=B8 
B9 18 19 jjmit  area=B9 
B10 22 16 jjmit  area=B10 
B11 23 24 jjmit  area=B11 
B12 26 27 jjmit  area=B12 
B13 29 30 jjmit  area=B13 
B14 32 31 jjmit  area=B14 
B15 33 34 jjmit  area=B15 
B16 36 37 jjmit  area=B16 
B17 32 38 jjmit  area=B17 
B18 30 39 jjmit  area=B18 
B19 40 41 jjmit  area=B19 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 25 pwl(0 0 5p IB5)
IB6 0 28 pwl(0 0 5p IB6)
IB7 0 35 pwl(0 0 5p IB7)
IB8 0 42 pwl(0 0 5p IB8)

LB1 3 1 LB1 
LB2 10 8 LB2 
LB3 14 7 LB3 
LB4 20 18 LB4 
LB5 25 23 LB5 
LB6 27 28 LB6 
LB7 35 33 LB7 
LB8 42 40 LB8 

L1 a 1 L1 
L2 1 4 L2 
L3 6 7 L3 
L4 b 8 L4 
L5 8 11 L5 
L6 7 13 L6 
L7 15 16 L7 
L8 clk 18 L8 
L9 18 21 L9 
L10 21 22 L10 
L11 16 23 L11 
L12 23 26 L12 
L13 27 29 L13 
L14 31 27 L14 
L15 21 33 L15 
L16 33 36 L16 
L17 36 32 L17 
L18 38 30 L18 
L19 30 40 L19 
L20 40 q L20 

LP1 2 0 LP1 
LP2 5 0 LP2 
LP4 9 0 LP4 
LP5 12 0 LP5 
LP8 17 0 LP8 
LP9 19 0 LP9 
LP11 24 0 LP11 
LP15 34 0 LP15 
LP16 37 0 LP16 
LP18 39 0 LP18 
LP19 41 0 LP19 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 4 106 RB3  
LRB3 106 6 LRB3 
RB4 8 108 RB4  
LRB4 108 0 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 11 113 RB6  
LRB6 113 13 LRB6 
RB7 7 115 RB7  
LRB7 115 15 LRB7 
RB8 16 116 RB8  
LRB8 116 0 LRB8 
RB9 18 118 RB9  
LRB9 118 0 LRB9 
RB10 22 122 RB10  
LRB10 122 16 LRB10 
RB11 23 123 RB11  
LRB11 123 0 LRB11 
RB12 26 126 RB12  
LRB12 126 27 LRB12 
RB13 29 129 RB13  
LRB13 129 30 LRB13 
RB14 32 131 RB14  
LRB14 131 31 LRB14 
RB15 33 133 RB15  
LRB15 133 0 LRB15 
RB16 36 136 RB16  
LRB16 136 0 LRB16 
RB17 32 138 RB17  
LRB17 138 38 LRB17 
RB18 30 130 RB18  
LRB18 130 0 LRB18 
RB19 40 140 RB19  
LRB19 140 0 LRB19 

.ends
