* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/07/29.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 29 July 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports a	b	q
.subckt THmitll_MERGE a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7'

.param B1=2.5
.param B2=3.01
.param B3=1.18
.param B4=2.5
.param B5=3.01
.param B6=1.18
.param B7=2.5

.param IB1=175u
.param IB2=175u
.param IB3=183u
.param IB4=175u

.param L1=2.0465p
.param L2=2.4953p
.param L3=0.9488p
.param L4=2.0465p
.param L5=2.4953p
.param L6=0.9488p
.param L7=3.6821p
.param L8=1.3761p

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB

.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP7=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 4 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 11 13 jjmit  area=B6 
B7 15 16 jjmit  area=B7 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 17 pwl(0 0 5p IB4)

LB1 3 1 LB1 
LB2 10 8 LB2 
LB3 14 7 LB3 
LB4 17 15 LB4 

L1 a 1 2.048E-012 
L2 1 4 2.485E-012 
L3 6 7 9.486E-013 
L4 b 8 2.059E-012 
L5 8 11 2.473E-012 
L6 7 13 9.53E-013 
L7 7 15 3.697E-012 
L8 15 q 1.377E-012 

LP1 2 0 4.88E-013 
LP2 5 0 3.854E-013 
LP4 9 0 4.857E-013 
LP5 12 0 3.834E-013 
LP7 16 0 3.61E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 4 106 RB3  
LRB3 106 6 LRB3 
RB4 8 108 RB4  
LRB4 108 0 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 11 113 RB6  
LRB6 113 13 LRB6 
RB7 15 115 RB7  
LRB7 115 0 LRB7 

.ends
