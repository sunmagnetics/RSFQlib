* Back-annotated simulation file written by InductEx v.6.0.4 on 3-6-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 3 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a q
.subckt LSmitll_PTLRX a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param LB=2p
.param Lptl=2p

.param B1=1
.param B2=1
.param B3=1

.param IB1=155u

.param L1=Lptl
.param L2=4.3p
.param L3=4.6p
.param L4=5p
.param L5=2.3p

.param LB1=LB
.param LP1=LP         
.param LP2=LP          
.param LP3=LP  

.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3   
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 3 8 jjmit area=B1
B2 4 10 jjmit area=B2
B3 5 12 jjmit area=B3

IB1 0 6 pwl(0 0 5p IB1)
LB1 6 7 3.274E-12
L1 a 3 1.499E-12
L2 3 7 4.327E-12
L3 7 4 4.63E-12
L4 4 5 4.962E-12
L5 5 q 2.298E-12

LP1 8 0 5.404E-13
LP2 10 0 6.269E-13
LP3 12 0 6.253E-13

RB1 3 9 RB1
RB2 4 11 RB2
RB3 5 13 RB3
LRB1 9 0 LRB1
LRB2 11 0 LRB2
LRB3 13 0 LRB3
.ends
