* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 26 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_ALWAYS0T_ASYNC_NOA_v3p0_base.cir
.endc

L1 1 q [L1]

* Ports
P1 q 0

PR1 1 0

.end