* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/07.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 4 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports 	a	b	clk	q
.subckt THmitll_OR2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=1.67
.param B3=1.48
.param B4=2.5
.param B5=1.67
.param B6=1.48
.param B7=2.27
.param B8=2.36
.param B9=1.76
.param B10=2.5
.param B11=1.44
.param B12=2.5

.param IB1=175u
.param IB2=175u
.param IB3=283u
.param IB4=158u
.param IB5=175u
.param IB6=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB

.param L1=1.6049p
.param L2=4.4173p
.param L3=0.7163p
.param L4=1.6049p
.param L5=4.4173p
.param L6=0.7163p
.param L7=3.2947p
.param L8=8.7190p
.param L9=2.1422p
.param L10=3.7843p
.param L11=3.9628p
.param L12=1.6906p

.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP8=LP
.param LP9=LP
.param LP10=LP
.param LP12=LP

.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10 
.param RB11=B0Rs/B11 
.param RB12=B0Rs/B12 

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 4 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 11 13 jjmit  area=B6 
B7 15 16 jjmit  area=B7 
B8 16 17 jjmit  area=B8 
B9 19 20 jjmit  area=B9 
B10 21 22 jjmit  area=B10 
B11 24 19 jjmit  area=B11 
B12 25 26 jjmit  area=B12 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)
IB6 0 27 pwl(0 0 5p IB6)

LB1 3 1 LB1 
LB2 10 8 LB2 
LB3 14 7 LB3 
LB4 18 16 LB4 
LB5 23 21 LB5 
LB6 27 25 LB6 

L1 a 1 1.592E-012 
L2 1 4 4.395E-012 
L3 6 7 7.134E-013 
L4 b 8 1.61E-012 
L5 8 11 4.378E-012 
L6 13 7 7.212E-013 
L7 7 15 3.29E-012 
L8 16 19 8.747E-012 
L9 clk 21 2.161E-012 
L10 21 24 3.766E-012 
L11 19 25 3.926E-012 
L12 25 q 1.675E-012 

LP1 2 0 4.683E-013 
LP2 5 0 4.125E-013 
LP4 9 0 3.472E-013 
LP5 12 0 4.43E-013 
LP8 17 0 4.666E-013 
LP9 20 0 4.384E-013 
LP10 22 0 3.63E-013 
LP12 26 0 4.421E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 4 106 RB3  
LRB3 106 6 LRB3 
RB4 8 108 RB4  
LRB4 108 0 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 11 113 RB6  
LRB6 113 13 LRB6 
RB7 15 115 RB7  
LRB7 115 16 LRB7 
RB8 16 116 RB8  
LRB8 116 0 LRB8 
RB9 19 119 RB9  
LRB9 119 0 LRB9 
RB10 21 121 RB10  
LRB10 121 0 LRB10 
RB11 24 124 RB11  
LRB11 124 19 LRB11 
RB12 25 125 RB12  
LRB12 125 0 LRB12 

.ends
