* Author: L. Schindler
* Version: 1.1.40
* Last modification date: 30 January 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

* Ports 			IN IN CLK OUT	
.subckt LSmitll_XORT a b clk q
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01=2.7984 
.param B01rx1=1.2124 
.param B01rx3=0.7236 
.param B02rx1=1.1586 
.param B02rx3=0.7720 
.param B02tx1=1.3695 
.param B03=1.9159 
.param B03rx1=0.8978 
.param B03rx3=0.8280 
.param B07=1.4857 
.param B08=0.9336 
.param B09=1.2859 
.param B10=1.6863 
.param IB01=8.9218e-05 
.param IB01rx1=0.000229789 
.param IB01rx3=0.000131858 
.param IB02tx1=6.64568e-05 
.param IB04=0.000134046 
.param IB05=0.000177629 
.param L01rx1=1.8604e-12 
.param L01rx3=1.8928e-12 
.param L02rx1=2.1529e-12 
.param L02rx3=2.2381e-12 
.param L03=2.2793e-12 
.param L03rx1=1.9729e-12 
.param L03rx3=2.0205e-12 
.param L03tx1=2.2261e-12 
.param L04rx1=2.3966e-12 
.param L04rx3=2.0178e-12 
.param L08=1.7515e-12 
.param L09=1.2620e-12 
.param L10=2.2246e-12 
.param L11=1.8033e-12 
.param L12=3.8658e-12 
.param L14=1.6354e-12 
.param LRB01=(RB01/Rsheet)*Lsheet
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01rx3=(RB01rx3/Rsheet)*Lsheet
.param LRB02rx1=(RB02rx1/Rsheet)*Lsheet
.param LRB02rx3=(RB02rx3/Rsheet)*Lsheet
.param LRB02tx1=(RB02tx1/Rsheet)*Lsheet
.param LRB03=(RB03/Rsheet)*Lsheet
.param LRB03rx1=(RB03rx1/Rsheet)*Lsheet
.param LRB03rx3=(RB03rx3/Rsheet)*Lsheet
.param LRB07=(RB07/Rsheet)*Lsheet
.param LRB08=(RB08/Rsheet)*Lsheet
.param LRB09=(RB09/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param RB01=B0Rs/B01
.param RB01rx1=B0Rs/B01rx1
.param RB01rx3=B0Rs/B01rx3
.param RB02rx1=B0Rs/B02rx1
.param RB02rx3=B0Rs/B02rx3
.param RB02tx1=B0Rs/B02tx1
.param RB03=B0Rs/B03
.param RB03rx1=B0Rs/B03rx1
.param RB03rx3=B0Rs/B03rx3
.param RB07=B0Rs/B07
.param RB08=B0Rs/B08
.param RB09=B0Rs/B09
.param RB10=B0Rs/B10
B01 10 49 78 jjmit area=B01
B01rx1 12 43 75 jjmit area=B01rx1
B01rx2 22 61 83 jjmit area=B01rx1
B01rx3 7 29 70 jjmit area=B01rx3
B02rx1 13 45 76 jjmit area=B02rx1
B02rx2 23 63 84 jjmit area=B02rx1
B02rx3 8 31 71 jjmit area=B02rx3
B02tx1 19 57 81 jjmit area=B02tx1
B03 10 11 74 jjmit area=B03
B03rx1 14 47 77 jjmit area=B03rx1
B03rx2 24 65 85 jjmit area=B03rx1
B03rx3 9 33 72 jjmit area=B03rx3
B04 20 67 86 jjmit area=B01
B06 20 21 82 jjmit area=B03
B07 16 17 79 jjmit area=B07
B08 18 55 80 jjmit area=B08
B09 5 6 69 jjmit area=B09
B10 5 35 73 jjmit area=B10
IB01 0 38 pwl(0 0 5p IB01)
IB01rx1 0 37 pwl(0 0 5p IB01rx1)
IB01rx2 0 53 pwl(0 0 5p IB01rx1)
IB01rx3 0 25 pwl(0 0 5p IB01rx3)
IB02 0 54 pwl(0 0 5p IB01)
IB02tx1 0 42 pwl(0 0 5p IB02tx1)
IB04 0 41 pwl(0 0 5p IB04)
IB05 0 26 pwl(0 0 5p IB05)
L01rx1 a 12 L01rx1
L01rx2 b 22 L01rx1
L01rx3 clk 7 L01rx3
L02rx1 12 39 L02rx1
L02rx2 22 59 L02rx1
L02rx3 7 27 L02rx3
L03 11 15 L03
L03rx1 39 13 L03rx1
L03rx2 59 23 L03rx1
L03rx3 27 8 L03rx3
L03tx1 19 52 L03tx1
L04rx1 13 14 L04rx1
L04rx2 23 24 L04rx1
L04rx3 8 9 L04rx3
L06 15 21 L03
L08 15 16 L08
L09 17 18 L09
L10 6 18 L10
L11 9 5 L11
L12 18 19 L12
L14 14 10 L14
L15 24 20 L14
LP01 49 0 2e-13
LP01rx1 43 0 2e-13
LP01rx2 61 0 2e-13
LP01rx3 29 0 2e-13
LP02rx1 45 0 2e-13
LP02rx2 63 0 2e-13
LP02rx3 31 0 2e-13
LP02tx1 57 0 2e-13
LP03 67 0 2e-13
LP03rx1 47 0 2e-13
LP03rx2 65 0 2e-13
LP03rx3 33 0 2e-13
LP05 55 0 2e-13
LP10 35 0 2e-13
LPR01 38 10 2e-13
LPR01rx1 37 39 2e-13
LPR01rx2 53 59 2e-13
LPR01rx3 25 27 2e-13
LPR02 54 20 2e-13
LPR02tx1 42 19 2e-13
LPR04 41 15 2e-13
LPR05 26 5 2e-13
LRB01 50 0 LRB01
LRB01rx1 44 0 LRB01rx1
LRB01rx2 62 0 LRB01rx1
LRB01rx3 30 0 LRB01rx3
LRB02rx1 46 0 LRB02rx1
LRB02rx2 64 0 LRB02rx1
LRB02rx3 32 0 LRB02rx3
LRB02tx1 58 0 LRB02tx1
LRB03 40 11 LRB03
LRB03rx1 48 0 LRB03rx1
LRB03rx2 66 0 LRB03rx1
LRB03rx3 34 0 LRB03rx3
LRB04 68 0 LRB01
LRB06 60 21 LRB03
LRB07 51 17 LRB07
LRB08 56 0 LRB08
LRB09 28 6 LRB09
LRB10 36 0 LRB10
RB01 10 50 RB01
RB01rx1 12 44 RB01rx1
RB01rx2 22 62 RB01rx1
RB01rx3 7 30 RB01rx3
RB02rx1 13 46 RB02rx1
RB02rx2 23 64 RB02rx1
RB02rx3 8 32 RB02rx3
RB02tx1 19 58 RB02tx1
RB03 10 40 RB03
RB03rx1 14 48 RB03rx1
RB03rx2 24 66 RB03rx1
RB03rx3 9 34 RB03rx3
RB04 20 68 RB01
RB06 20 60 RB03
RB07 16 51 RB07
RB08 18 56 RB08
RB09 5 28 RB09
RB10 5 36 RB10
RINStx1 52 q 1.36
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.ends LSmitll_XORT
