* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===
*$Ports  a b clk q
.subckt LSMITLL_AND2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param B2=IC/1.4
.param B3=IC
.param B4=IC/1.4
.param B5=IC
.param B6=IC/1.4
.param B7=B1
.param B8=B2
.param B9=B3
.param B10=B4
.param B11=B5
.param B12=B6
.param B13=IC
.param B14=IC
.param B15=IC
.param IB1=BiasCoef*Ic0*B1
.param IB2=BiasCoef*Ic0*B3
.param IB3=IB1
.param IB4=IB2
.param IB5=BiasCoef*Ic0*B13
.param IB6=BiasCoef*Ic0*B14
.param IB7=BiasCoef*Ic0*B15
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(B3*Ic0)
.param L4=1p
.param L5=Phi0/(2*B5*Ic0)
.param L6=L1
.param L7=L2
.param L8=L3
.param L9=L4
.param L10=L5
.param L11=Phi0/(4*IC*Ic0)
.param L12=Phi0/(2*B13*Ic0)
.param L13=1p
.param L14=1p
.param L15=Phi0/(4*IC*Ic0)
.param LP1=LP
.param LP3=LP
.param LP5=LP
.param LP7=LP
.param LP9=LP
.param LP11=LP
.param LP13=LP
.param LP14=LP
.param LP15=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet
B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 8 11 jjmit area=B5
B6 12 13 jjmit area=B6
B7 14 15 jjmit area=B7
B8 17 18 jjmit area=B8
B9 18 19 jjmit area=B9
B10 21 22 jjmit area=B10
B11 21 23 jjmit area=B11
B12 24 13 jjmit area=B12
B13 25 26 jjmit area=B13
B14 31 32 jjmit area=B14
B15 28 29 jjmit area=B15
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 27 pwl(0 0 5p IB5)
IB6 0 33 pwl(0 0 5p IB6)
IB7 0 30 pwl(0 0 5p IB7)
LB1 3 1 LB1
LB2 7 5 LB2
LB3 16 14 LB3
LB4 20 18 LB4
LB5 27 25 LB5
LB6 30 28 LB6
LB7 33 31 LB7
LP1 2 0 LP1
LP3 6 0 LP3
LP5 11 0 LP5
LP7 15 0 LP7
LP9 19 0 LP9
LP11 23 0 LP11
LP13 26 0 LP13
LP14 32 0 LP14
LP15 29 0 LP15
L1 a 1 L1
L2 1 4 L2
L3 5 8 L3
L4 9 10 L4
L5 8 12 L5
L6 b 14 L6
L7 14 17 L7
L8 18 21 L8
L9 22 10 L9
L10 21 24 L10
L11 clk 25 L11
L12 25 31 L12
L13 31 10 L13
L14 13 28 L14
L15 28 q L15
RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 5 105 RB3
LRB3 105 0 LRB3
RB4 8 109 RB4
LRB4 109 9 LRB4
RB5 8 108 RB5
LRB5 108 0 LRB5
RB6 12 112 RB6
LRB6 112 13 LRB6
RB7 14 114 RB7
LRB7 114 0 LRB7
RB8 17 117 RB8
LRB8 117 18 LRB8
RB9 18 118 RB9
LRB9 118 0 LRB9
RB10 21 122 RB10
LRB10 122 22 LRB10
RB11 21 121 RB11
LRB11 121 0 LRB11
RB12 24 124 RB12
LRB12 124 13 LRB12
RB13 25 125 RB13
LRB13 125 0 LRB13
RB14 31 131 RB14
LRB14 131 0 LRB14
RB15 28 128 RB15
LRB15 128 0 LRB15
.ends
* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 11
b1   1  2  jjmitll100 area=2.25
b2   3  4  jjmitll100 area=2.25
b3   5  6  jjmitll100 area=2.5
ib1  0  2  pwl(0 0 5p 275ua)
ib2  0  5  pwl(0 0 5p 175ua)
l1   8  7  1p
l2   7  0  3.9p
l3   7  1  0.6p
l4   2  3  1.1p
l5   3  5  4.5p
l6   5  11 2p
lp2  4  0  0.2p
lp3  6  0  0.2p
lrb1 9  2  1p
lrb2 10 4  1p
lrb3 12 6  1p
rb1  1  9  4.31
rb2  3  10 4.31
rb3  5  12 3.88
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.2p
.param ic=2.5
.param icreceive=2.5
.param ictrans=2.5
.param lptl=2p
.param lb=2p
.param biascoef=0.7
.param b1=ic
.param b2=ic
.param rb1=b0rs/b1
.param rb2=b0rs/b2
.param lrb1=(rb1/rsheet)*lsheet
.param lrb2=(rb2/rsheet)*lsheet
.param l1=lptl
.param l2=phi0/(4*b1*ic0)
.param l3=phi0/(4*b1*ic0)
.param l4=lptl
.param ib1=biascoef*ic0*(b1+b2)
b1  3 7 jjmit  area=b1
b2 4 9 jjmit  area=b2
ib1 0 5 pwl(0 0 5p ib1)
l1 a 3 l1
l2 3 6 l2
l3 6 4 l3
l4 4 q l4
lb1 5 6 lb
lp1 7 0 lp
lp2 9 0 lp
lrb1 3 8 lrb1
lrb2 4 10 lrb2
rb1 8 0 rb1
rb2 10 0 rb2
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.2p
.param ic=2.5
.param icreceive=2.5
.param ictrans=2.5
.param lptl=2p
.param lb=2p
.param biascoef=0.7
.param b1=ic
.param b2=ic
.param rb1=b0rs/b1
.param rb2=b0rs/b2
.param lrb1=(rb1/rsheet)*lsheet
.param lrb2=(rb2/rsheet)*lsheet
.param l1=lptl
.param l2=phi0/(4*b1*ic0)
.param l3=phi0/(4*b1*ic0)
.param l4=lptl
.param ib1=biascoef*ic0*(b1+b2)
b1  3 7 jjmit  area=b1
b2 4 9 jjmit  area=b2
ib1 0 5 pwl(0 0 5p ib1)
l1 a 3 l1
l2 3 6 l2
l3 6 4 l3
l4 4 q l4
lb1 5 6 lb
lp1 7 0 lp
lp2 9 0 lp
lrb1 3 8 lrb1
lrb2 4 10 lrb2
rb1 8 0 rb1
rb2 10 0 rb2
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  1
r1 1 0 2
.ENDS SINKCELL
* ===== MAIN =====
I_a 0 1001 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa SOURCECELL 1001 1002
XLOADINa LOADINCELL 1002 a
I_b 0 1004 pwl(0 0 350p 0 353p 600u 356p 0 450p 0 453p 600u 456p 0 480p 0 483p 600u 486p 0 560p 0 563p 600u 566p 0 580p 0 583p 600u 586p 0 660p 0 663p 600u 666p 0 740p 0 743p 600u 746p 0)
XSOURCEINb SOURCECELL 1004 1005
XLOADINb LOADINCELL 1005 b
I_clk 0 1007 pulse(0 600u 20p 2p 2p 1p 100p)
XSOURCEINclk SOURCECELL 1007 1008
XLOADINclk LOADINCELL 1008 clk
XLOADOUTq LOADOUTCELL q 10011
XSINKOUTq SINKCELL 10011
XDUT lsmitll_and2 a b clk q
.tran 0.025p 1000p 0
.print i(L1.XDUT) p(B1.XDUT) i(L6.XDUT) p(B7.XDUT) i(L11.XDUT) p(B13.XDUT) p(B15.XDUT) p(B1.XLOADOUTq)
.end
