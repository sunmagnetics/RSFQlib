* Back-annotated simulation file written by InductEx v.6.0.4 on 27-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 26 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a q
.subckt LSmitll_PTLRX_SFQDC a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=2p
.param LP=0.2p

.param B1=1
.param B2=1
.param B3=1
.param B4=3.25
.param B5=1.50
.param B6=1.75
.param B7=2.00
.param B8=3.00
.param B9=1.50
.param B10=1.50
.param B11=2.00

.param IB1=155u
.param IB2=280u
.param IB3=150u
.param IB4=220u
.param IB5=80u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet

.param R1=5.74


B1 2 3 jjmit area=B1
B2 6 7 jjmit area=B2
B3 8 9 jjmit area=B3
B4 10 11 jjmit area=B4
B5 13 14 jjmit area=B5
B6 15 16 jjmit area=B6
B7 19 20 jjmit area=B7
B8 20 21 jjmit area=B8
B9 23 24 jjmit area=B9
B10 26 27 jjmit area=B10
B11 30 31 jjmit area=B11

LP1 3 0 5.068E-13
LP2 7 0 6.182E-13
LP3 9 0 6.097E-13
LP4 11 0 4.785E-13
LP6 16 0 4.984E-13
LP8 21 0 4.692E-13
LP10 27 0 5.018E-13
LP11 31 0 5.645E-13

IB1 0 5 pwl(0 0 5p IB1)
IB2 0 12 pwl(0 0 5p IB2)
IB3 0 17 pwl(0 0 5p IB3)
IB4 0 25 pwl(0 0 5p IB4)
IB5 0 29 pwl(0 0 5p IB5)

LB1 4 5 1.284E-12
LB2 10 12 3.934E-12
LB3 15 17 1.916E-12
LB4 24 25 5.378E-12
LB5 28 29 3.797E-12

L1 a 2 1.524E-12
L2 2 4 4.301E-12
L3 4 6 4.612E-12
L4 6 8 5.035E-12
L5 8 10 3.791E-12
L6 10 13 8.316E-13
L7 14 15 1.167E-12
L9 15 18 5.964E-12
L10 13 19 1.104E-12
L11 20 18 3.24E-12
L12 18 22 8.87E-13
L14 18 23 5.769E-13
L15 24 26 9.383E-13
L16 26 28 3.701E-12
L17 28 30 2.06E-12
L18 30 q 4.08E-12

R1 22 0 R1

RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 6 106 RB2
LRB2 106 0 LRB2
RB3 8 108 RB3
LRB3 108 0 LRB3
RB4 10 110 RB4
LRB4 110 0 LRB4
RB5 13 113 RB5
LRB5 113 14 LRB5
RB6 15 115 RB6
LRB6 115 0 LRB6
RB7 19 119 RB7
LRB7 119 20 LRB7
RB8 20 120 RB8
LRB8 120 0 LRB8
RB9 23 123 RB9
LRB9 123 24 LRB9
RB10 26 126 RB10
LRB10 126 0 LRB10
RB11 30 130 RB11
LRB11 130 0 LRB11

.ends
