* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

*$Ports 			  a clk q
.subckt LSMITLL_DFFT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param ICreceive=2.0
.param ICtrans=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param RD=1.36
.param B1=ICreceive
.param B2=IC
.param B3=IC/1.4
.param B4=IC
.param B5=IC
.param B6=ICreceive
.param B7=IC
.param B8=IC/1.4
.param B9=IC
.param B10=ICtrans
.param IB1=BiasCoef*(B1*Ic0+B2*Ic0)
.param IB2=IC*Ic0
.param IB3=BiasCoef*(B6*Ic0+B7*Ic0)
.param IB4=BiasCoef*(B9*Ic0+B10*Ic0)
.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))/2
.param L3=(Phi0/(2*B1*Ic0))/2
.param L4=Phi0/(2*B2*Ic0)
.param L5=Phi0/(B4*Ic0)
.param L6=Lptl
.param L7=(Phi0/(2*B6*Ic0))/2
.param L8=(Phi0/(2*B6*Ic0))/2
.param L9=Phi0/(2*B7*Ic0)
.param L10=Phi0/(2*B5*Ic0)
.param L11=(Phi0/(2*B9*Ic0))/2
.param L12=(Phi0/(2*B9*Ic0))/2
.param L13=Lptl
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP9=LP
.param LP10=LP
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
IB1 0 5 pwl(0 0 5p IB1)
IB2 0 11 pwl(0 0 5p IB2)
IB3 0 18 pwl(0 0 5p IB3)
IB4 0 25 pwl(0 0 5p IB4)
B1 2 3 jjmit area=B1
B2 6 7 jjmit area=B2
B3 8 9 jjmit area=B3
B4 9 10 jjmit area=B4
B5 12 13 jjmit area=B5
B6 15 16 jjmit area=B6
B7 19 20 jjmit area=B7
B8 21 12 jjmit area=B8
B9 22 23 jjmit area=B9
B10 26 27 jjmit area=B10
L1 a 2 L1
L2 2 4 L2
L3 4 6 L3
L4 6 8 L4
L5 9 12 L5
L6 clk 15 L6
L7 15 17 L7
L8 17 19 L8
L9 19 21 L9
L10 12 22 L10
L11 22 24 L11
L12 24 26 L12
L13 26 28 L13
LP1 3 0 LP1
LP2 7 0 LP2
LP4 10 0 LP4
LP5 13 0 LP5
LP6 16 0 LP6
LP7 20 0 LP7
LP9 23 0 LP9
LP10 27 0 LP10
LB1 4 5 LB1
LB2 9 11 LB2
LB3 17 18 LB3
LB4 24 25 LB4
RB1 2 102 RB1
RB2 6 106 RB2
RB3 8 108 RB3
RB4 9 109 RB4
RB5 12 112 RB5
RB6 15 115 RB6
RB7 19 119 RB7
RB8 21 121 RB8
RB9 22 122 RB9
RB10 26 126 RB10
LRB1 102 0 LRB1
LRB2 106 0 LRB2
LRB3 108 9 LRB3
LRB4 109 0 LRB4
LRB5 112 0 LRB5
LRB6 115 0 LRB6
LRB7 119 0 LRB7
LRB8 121 12 LRB8
LRB9 122 0 LRB9
LRB10 126 0 LRB10
RD 28 q RD
.ends