* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/09.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 14 April 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	q
.subckt THmitll_DCSFQ-PTLTX a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=0.9*Ic
.param B2=0.9*Ic
.param B3=IC
.param B4=ICtrans

.param IB1=(11/9)*Ic0*B2
.param IB2=BiasCoef*Ic0*(B3+B4)

.param LB1=LB
.param LB2=LB

.param LP2=LP
.param LP3=LP
.param LP4=LP

.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=Phi0/(2*B2*Ic0)
.param L6=Phi0/(4*B3*Ic0)
.param L7=Phi0/(4*B3*Ic0)
.param L8=Lptl

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP

B1 2 3 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 11 12 jjmit  area=B4 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)

LB1 4 3 3.12E-012 
LB2 10 9 8.782E-013 

LP2 6 0 5.209E-013 
LP3 8 0 5.058E-013 
LP4 12 0 4.053E-013 

L1 a 1 1.322E-012 
L2 1 0 3.879E-012 
L3 1 2 6.03E-013 
L4 3 5 1.104E-012 
L5 5 7 4.572E-012 
L6 7 9 2.078E-012 
L7 9 11 2.073E-012 
L8 11 13 8.436E-013 

RD 13 q RD  

RB1 2 102 RB1  
LRB1 102 3 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 11 111 RB4  
LRB4 111 0 LRB4 

.ends
