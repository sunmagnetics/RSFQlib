* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===
* Back-annotated simulation file written by InductEx v.6.0.4 on 27-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 8 June 2021
* Last modification by: L. Schindler
* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University
* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:
* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.
* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.
* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za
*$Ports 			  a clk q
.subckt LSMITLL_DFFT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param ICreceive=2.0
.param ICtrans=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param RD=1.36

.param B1=1.62
.param B2=1.89
.param B3=1.72
.param B4=2.32
.param B5=2.12
.param B6=1.62
.param B7=1.98
.param B8=1.71
.param B9=2.12
.param B10=2.5

.param IB1=276u
.param IB2=235u
.param IB3=284u
.param IB4=312u

.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))/2
.param L3=(Phi0/(2*B1*Ic0))/2
.param L4=Phi0/(2*B2*Ic0)
.param L5=Phi0/(B4*Ic0)
.param L6=Lptl
.param L7=(Phi0/(2*B6*Ic0))/2
.param L8=(Phi0/(2*B6*Ic0))/2
.param L9=Phi0/(2*B7*Ic0)
.param L10=Phi0/(2*B5*Ic0)
.param L11=(Phi0/(2*B9*Ic0))/2
.param L12=(Phi0/(2*B9*Ic0))/2
.param L13=Lptl
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP9=LP
.param LP10=LP
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
IB1 0 5 pwl(0 0 5p IB1)
IB2 0 11 pwl(0 0 5p IB2)
IB3 0 18 pwl(0 0 5p IB3)
IB4 0 25 pwl(0 0 5p IB4)
B1 2 3 jjmit area=B1
B2 6 7 jjmit area=B2
B3 8 9 jjmit area=B3
B4 9 10 jjmit area=B4
B5 12 13 jjmit area=B5
B6 15 16 jjmit area=B6
B7 19 20 jjmit area=B7
B8 21 12 jjmit area=B8
B9 22 23 jjmit area=B9
B10 26 27 jjmit area=B10
L1 a 2 1.587E-12
L2 2 4 3.253E-12
L3 4 6 3.304E-12
L4 6 8 3.979E-12
L5 9 12 7.521E-12
L6 clk 15 1.6E-12
L7 15 17 3.042E-12
L8 17 19 3.045E-12
L9 19 21 4.21E-12
L10 12 22 4.022E-12
L11 22 24 2.164E-12
L12 24 26 2.183E-12
L13 26 28 2.536E-12
LP1 3 0 5.021E-13
LP2 7 0 5.102E-13
LP4 10 0 5.275E-13
LP5 13 0 5.37E-13
LP6 16 0 5.005E-13
LP7 20 0 5.161E-13
LP9 23 0 5.212E-13
LP10 27 0 5.039E-13
LB1 4 5 3.559E-12
LB2 9 11 2.45E-12
LB3 17 18 2.72E-12
LB4 24 25 1.988E-12
RB1 2 102 RB1
RB2 6 106 RB2
RB3 8 108 RB3
RB4 9 109 RB4
RB5 12 112 RB5
RB6 15 115 RB6
RB7 19 119 RB7
RB8 21 121 RB8
RB9 22 122 RB9
RB10 26 126 RB10
LRB1 102 0 LRB1
LRB2 106 0 LRB2
LRB3 108 9 LRB3
LRB4 109 0 LRB4
LRB5 112 0 LRB5
LRB6 115 0 LRB6
LRB7 119 0 LRB7
LRB8 121 12 LRB8
LRB9 122 0 LRB9
LRB10 126 0 LRB10
RD 28 q RD
.ends
* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 22
b1    1  2  jjmitll100 area=2.25
b2    3  4  jjmitll100 area=2.25
b3    5  6  jjmitll100 area=2.5
ib1   0  2  pwl(0 0 5p 275ua)
ib2   0  5  pwl(0 0 5p 175ua)
l1    8  7  1p
l2    7  0  3.9p
l3    7  1  0.6p
l4    2  3  1.1p
l5    3  5  4.5p
l6    5  11 2p
lp2   4  0  0.2p
lp3   6  0  0.2p
lrb1  9  2  1p
lrb2  10 4  1p
lrb3  12 6  1p
rb1   1  9  4.31
rb2   3  10 4.31
rb3   5  12 3.88
b01   23 27 jjmitll100 area=2
b02   24 26 jjmitll100 area=1.62
ib01  0  30 pwl(0      0 5p 0.00023)
ib02  0  31 pwl(0      0 5p 8.2e-005)
l01   11 23 2.5e-012
l02   23 24 3.3e-012
l03   24 25 3.5e-013
lp01  0  27 5e-014
lp02  0  26 1.2e-013
lpr01 23 30 2e-013
lpr02 24 31 1.3e-012
lrb01 27 28 1e-012
lrb02 26 29 1e-012
rb01  28 23 4.85
rb02  29 24 6.3
rins  25 22 1.36
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
tload 2 0 5 0 lossless z0=5 td=10p
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
tload 2 0 5 0 lossless z0=5 td=50p
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  2
b1    1  9  jjmitll100     area=1
b2    4  8  jjmitll100     area=1
b3    5  7  jjmitll100     area=1
ib1   0  10 pwl(0      0 5p 145u)
l1    2  1  0.2p
l2    1  3  4.3p
l3    3  4  4.6p
l4    4  5  6.0p
l5    5  6  1.3p
lp1   0  9  0.34p
lp2   0  8  0.06p
lp3   0  7  0.03p
lpr1  3  10 0.2p
lrb1  9  11 0.5p
lrb2  8  12 1p
lrb3  7  13 1p
rb1   11 1  15.4
rb2   12 4  11.3
rb3   13 5  11.3
rsink 6  0  2
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160ohm, rn=16ohm, icrit=0.1ma)
.ENDS SINKCELL
* ===== MAIN =====
I_a 0 1 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa SOURCECELL 1 2
XLOADINa LOADINCELL 2 3
I_clk 0 4 pulse(0 600u 20p 2p 2p 1p 100p)
XSOURCEINclk SOURCECELL 4 5
XLOADINclk LOADINCELL 5 6
XLOADOUTq LOADOUTCELL 7 8
XSINKOUTq SINKCELL 8
XDUT lsmitll_dfft 3 6 7
.tran 0.025p 1000p 0
.print i(L1.XDUT) p(B1.XDUT) i(L6.XDUT) p(B6.XDUT) i(L13.XDUT) p(B10.XDUT)
.end
