* Author: L. Schindler
* Version: 2.1
* Last modification date: 28 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$ports a b clk q
.subckt LSMITLL_OR2T a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param Lptl=2p
.param LB=2p
.param RD=1.36

.param B1=1.17
.param B2=1.95
.param B3=1.31
.param B4=1.17
.param B5=1.95
.param B6=1.31
.param B7=2.20
.param B8=1.72
.param B9=0.81
.param B10=0.75
.param B11=0.63
.param B12=1.40
.param B13=1.62
.param B14=1.9

.param IB1=141u
.param IB2=141u
.param IB3=328u
.param IB4=81u
.param IB5=98u
.param IB6=81u
.param IB7=177u

.param L1=Lptl
.param L2=2.0822p
.param L3=2.6809p
.param L4=1.3486p
.param L5=Lptl
.param L6=2.0822p
.param L7=2.6809p
.param L8=1.3486p	
.param L10=1.8890p
.param L12=5.4916p
.param L13=Lptl
.param L14=3.3652p
.param L15=4.0267p	
.param L16=0.7p
.param L17=1.5727p
.param L18=2.0776p
.param L19=0.885p
.param L20=4.2904p	
.param L21=Lptl

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP8=LP
.param LP9=LP
.param LP10=LP
.param LP12=LP
.param LP13=LP
.param LP14=LP

.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11   
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
.param LRB12=(RB12/Rsheet)*Lsheet+LP
.param LRB13=(RB13/Rsheet)*Lsheet+LP
.param LRB14=(RB14/Rsheet)*Lsheet+LP

B1 2 3  	jjmit area=B1
B2 6 7  	jjmit area=B2
B3 6 8		jjmit area=B3
B4 11 12	jjmit area=B4
B5 15 16	jjmit area=B5
B6 15 43	jjmit area=B6
B7 19 22	jjmit area=B7
B8 22 21	jjmit area=B8
B9 26 27	jjmit area=B9
B10 30 31	jjmit area=B10
B11 32 24	jjmit area=B11
B12 33 34	jjmit area=B12
B13 37 38	jjmit area=B13
B14 39 41	jjmit area=B14

IB1 0 5  pwl(0 0 5p IB1)
IB2 0 14 pwl(0 0 5p IB2)
IB3 0 18 pwl(0 0 5p IB3)
IB4 0 23 pwl(0 0 5p IB4)
IB5 0 29 pwl(0 0 5p IB5)
IB6 0 36 pwl(0 0 5p IB6)
IB7 0 40 pwl(0 0 5p IB7)

L1 a 2 L1		
L2 2 4 L2	
L3 4 6 L3	
L4 8 9 L4	
L5 b 11 L5			
L6 11 13 L6	
L7 13 15 L7		
L8 43 9 L8		
L10 9 19 L10	
L12 22 24 L12	
L13 clk 26 L13		
L14 26 28 L14	
L15 28 30 L15	
L16 30 32 L16	
L17 24 33 L17	
L18 33 35 L18	
L19 35 37 L19	
L20 37 39 L20	
L21 39 42 L21	
RD 42 q RD

LB1 4 5 LB1
LB2 13 14 LB2
LB3 9 18 LB3
LB4 22 23 LB4
LB5 28 29 LB5
LB6 35 36 LB6
LB7 39 40 LB7
LP1 3 0 LP1
LP2 7 0 LP2
LP4 12 0 LP4
LP5 16 0 LP5
LP8 21 0 LP8
LP9 27 0 LP9
LP10 31 0 LP10
LP12 34 0 LP12
LP13 38 0 LP13
LP14 41 0 LP14

RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 6 106 RB2
LRB2 106 0 LRB2
RB3 6 108 RB3
LRB3 108 8 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
RB5 15 115 RB5
LRB5 115 0 LRB5
RB6 15 143 RB6
LRB6 143 43 LRB6
RB7 19 119 RB7
LRB7 119 22 LRB7
RB8 22 122 RB8
LRB8 122 0 LRB8
RB9 26 126 RB9
LRB9 126 0 LRB9
RB10 30 130 RB10
LRB10 130 0 LRB10
RB11 32 132 RB11
LRB11 132 24 LRB11
RB12 33 133 RB12
LRB12 133 0 LRB12
RB13 37 137 RB13
LRB13 137 0 LRB13
RB14 39 139 RB14
LRB14 139 0 LRB14
.ends
