* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 16 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_DFFT_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 [L1]
L2 1 3 2.8908p [L2]
L3 3 5 3.6865p [L3]
L4 5 7 4.7771p [L4]
L5 8 11 9.5023p [L5]
L6 clk 12 [L6]
L7 12 14 2.2014p [L7] 
L8 14 16 5.6199p [L8]
L9 16 18 5.3129p [L9]
L10 11 20 4.5588p [L10]
L11 20 q [L11]

LP1 2 0 [LP1] 
LP2 6 0 [LP2]
LP4 9 0 [LP4]
LP5 13 0 [LP5]
LP6 17 0 [LP6]
LP8 19 0 [LP8]
LP9 21 0 [LP9]

LB1 4 3 [LB1]
LB2 10 8 [LB2]
LB3 14 15 [LB3]
LB4 20 22 [LB4]

* Ports
P1 a 0
P2 clk 0
P3 q 0

PB1 4 0
PB2 10 0
PB3 15 0
PB4 22 0

J1 1 2		160u
J2 5 6 		182u
J3 7 8		136u
J4 8 9		207u
J5 12 13	160u
J6 16 17	127u
J7 18 11	128u
J8 11 19	189u
J9 20 21	250u

.end
