* Back-annotated simulation file written by InductEx v.6.0.4 on 2-6-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 2 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a q
.subckt LSmitll_DCSFQ_PTLTX a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LB=0.2p
.param LP=0.2p
.param B1=2.25
.param B2=2.25
.param B3=2.5
.param B4=2
.param B5=1.62
.param IB1=275u
.param IB2=175u
.param IB3=230u
.param IB4=82u
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=4.5p
.param L7=3.3p
.param L8=0.35p
.param RD=1.36
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 6 7 jjmit area=B2
B3 9 10 jjmit area=B3
B4 13 14 jjmit area=B4
B5 17 18 jjmit area=B5
IB1 0 5 pwl(0 0 5p IB1)
IB2 0 12 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
LB1 5 3 3.122E-12
LB2 12 9 2.229E-12
LB3 16 13 6.294E-13
LB4 20 17 2.139E-12
L1 a 1 1.293E-12
L2 1 0 3.9E-12
L3 1 2 5.991E-13
L4 3 6 1.088E-12
L5 6 9 4.514E-12
L6 9 13 4.542E-12
L7 13 17 3.272E-12
L8 17 21 1.009E-12
LP2 7 0 5.238E-13
LP3 10 0 5.263E-13
LP4 14 0 4.571E-13
LP5 18 0 4.763E-13
LRB1 2 4 LRB1
LRB2 8 0 LRB2
LRB3 11 0 LRB3
LRB4 15 0 LRB4
LRB5 19 0 LRB5
RB1 4 3 RB1
RB2 6 8 RB2
RB3 9 11 RB3
RB4 13 15 RB4
RB5 17 19 RB5
RD 21 q RD
.ends
