* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===
* Back-annotated simulation file written by InductEx v.6.0.4 on 27-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 27 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$ports				   a b q
.subckt LSmitll_MERGET a b q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.70
.param RD=1.36

.param B1=1.6
.param B2=1.54
.param B3=0.95
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=1.16
.param B8=2.5
.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)*(B7/(B2+B7))
.param L4=L1
.param L5=L2
.param L6=L3
.param L7=Phi0/(2*B2*Ic0)*(B2/(B2+B7))
.param L8=(Phi0/(2*B7*Ic0))*(B8/(B7+B8))
.param L9=(Phi0/(2*B7*Ic0))*(B7/(B7+B8))
.param L10=Lptl
.param IB1=148u
.param IB2=148u
.param IB3=241u
.param IB4=176u
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet

L1 a 1 1.439E-12
L2 1 4 6.953E-12
L3 4 6 1.156E-12
L4 b 8 1.462E-12
L5 8 11 6.998E-12
L6 11 13 1.166E-12
L7 7 15 3.436E-12
L8 15 19 2.713E-12
L9 17 19 2.713E-12
L10 19 21 7.598E-13
RD 21 q RD
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 6 7 jjmit area=B3
B4 8 9 jjmit area=B4
B5 11 12 jjmit area=B5
B6 13 7 jjmit area=B6
B7 15 16 jjmit area=B7
B8 19 20 jjmit area=B8
LP1 2 0 4.853E-13
LP2 5 0 5.381E-13
LP4 9 0 4.789E-13
LP5 12 0 5.351E-13
LP7 16 9 5.981E-13
LP8 20 0 3.813E-13
RB1 1 101 RB1
RB2 4 104 RB2
RB3 6 106 RB3
RB4 8 108 RB4
RB5 11 111 RB5
RB6 13 113 RB6
RB7 15 115 RB7
RB8 19 119 RB8
LRB1 101 0 LRB1
LRB2 104 0 LRB2
LRB3 106 7 LRB3
LRB4 108 0 LRB4
LRB5 111 0 LRB5
LRB6 113 7 LRB6
LRB7 115 0 LRB7
LRB8 119 0 LRB8
LB1 1 3 2.952E-12
LB2 8 10 2.928E-12
LB3 7 14 2.643E-12
LB4 17 18 1.428E-12
.ends

* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 22
b1    1  2  jjmitll100 area=2.25
b2    3  4  jjmitll100 area=2.25
b3    5  6  jjmitll100 area=2.5
ib1   0  2  pwl(0 0 5p 275ua)
ib2   0  5  pwl(0 0 5p 175ua)
l1    8  7  1p
l2    7  0  3.9p
l3    7  1  0.6p
l4    2  3  1.1p
l5    3  5  4.5p
l6    5  11 2p
lp2   4  0  0.2p
lp3   6  0  0.2p
lrb1  9  2  1p
lrb2  10 4  1p
lrb3  12 6  1p
rb1   1  9  4.31
rb2   3  10 4.31
rb3   5  12 3.88
b01   23 27 jjmitll100 area=2
b02   24 26 jjmitll100 area=1.62
ib01  0  30 pwl(0      0 5p 0.00023)
ib02  0  31 pwl(0      0 5p 8.2e-005)
l01   11 23 2.5e-012
l02   23 24 3.3e-012
l03   24 25 3.5e-013
lp01  0  27 5e-014
lp02  0  26 1.2e-013
lpr01 23 30 2e-013
lpr02 24 31 1.3e-012
lrb01 27 28 1e-012
lrb02 26 29 1e-012
rb01  28 23 4.85
rb02  29 24 6.3
rins  25 22 1.36
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
tload 2 0 5 0 lossless z0=5 td=10p
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
tload 2 0 5 0 lossless z0=5 td=50p
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  2
b1    1  9  jjmitll100     area=1
b2    4  8  jjmitll100     area=1
b3    5  7  jjmitll100     area=1
ib1   0  10 pwl(0      0 5p 145u)
l1    2  1  0.2p
l2    1  3  4.3p
l3    3  4  4.6p
l4    4  5  6.0p
l5    5  6  1.3p
lp1   0  9  0.34p
lp2   0  8  0.06p
lp3   0  7  0.03p
lpr1  3  10 0.2p
lrb1  9  11 0.5p
lrb2  8  12 1p
lrb3  7  13 1p
rb1   11 1  15.4
rb2   12 4  11.3
rb3   13 5  11.3
rsink 6  0  2
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160ohm, rn=16ohm, icrit=0.1ma)
.ENDS SINKCELL
* ===== MAIN =====
I_a 0 1 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa SOURCECELL 1 2
XLOADINa LOADINCELL 2 3
I_b 0 4 pwl(0 0 350p 0 353p 600u 356p 0 450p 0 453p 600u 456p 0 480p 0 483p 600u 486p 0 560p 0 563p 600u 566p 0 580p 0 583p 600u 586p 0 660p 0 663p 600u 666p 0 740p 0 743p 600u 746p 0)
XSOURCEINb SOURCECELL 4 5
XLOADINb LOADINCELL 5 6
XLOADOUTq LOADOUTCELL 7 8
XSINKOUTq SINKCELL 8
XDUT lsmitll_merget 3 6 7
.tran 0.025p 1000p 0
.print i(L1.XDUT) p(B1.XDUT) i(L4.XDUT) p(B4.XDUT) i(L10.XDUT) p(B8.XDUT)
.end
