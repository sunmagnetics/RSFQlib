* Back-annotated simulation file written by InductEx v.6.0.4 on 3-6-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 24 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a q
.subckt LSmitll_PTLTX a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param LB=2p
.param Lptl=2p
.param RD=1.36

.param B1=2
.param B2=1.62

.param IB1=230u        
.param IB2=82u     

.param L1=2.5p            
.param L2=3.3p        
.param L3=Lptl
    
.param LB1=LB           
.param LB2=LB   
.param LP1=LP         
.param LP2=LP 
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2   
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet

B1 3 8 jjmit area=B1
B2 4 10 jjmit area=B2
IB1 0 5 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
LB1 5 3 2.86E-12
LB2 6 4 3.424E-12
L1 a 3 2.256E-12
L2 3 4 3.32E-12
L3 4 7 1.026E-12
RD 7 q RD
LP1 8 0 5.122E-13
LP2 10 0 4.727E-13
RB1 3 9 RB1
RB2 4 11 RB2
LRB1 9 0 LRB1
LRB2 11 0 LRB2
.ends
