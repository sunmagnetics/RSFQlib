* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 28 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_XOR_v3p0_optimised.cir
.endc

*Inductors
L1 a 1 1.5740p [L1]
L2 1 4 3.1407p [L2]
L3 6 7 4.7381p [L3]
L4 b 8 1.5740p [L4]
L5 8 11 3.1407p [L5]
L6 7 13 4.7381p [L6]
L7 15 16 4.7751p [L7]
L8 clk 18 1.1983p [L8]
L9 18 21 3.2191p [L9]
L10 16 22 3.7711p [L10]
L11 22 q 1.4703p [L11]

LP1 2 0 [LP1] 
LP2 5 0 [LP2] 
LP4 9 0 [LP4] 
LP5 12 0 [LP5] 
LP8 17 0 [LP8] 
LP9 19 0 [LP9] 
LP11 23 0 [LP11] 

LB1 3 1 [LB1] 
LB2 10 8 [LB2] 
LB3 14 7 [LB3] 
LB4 20 18 [LB4]
LB5 24 22 [LB5] 

*Ports
P1 a 0
P2 b 0
P3 clk 0
P4 q 0

PB1 3 0
PB2 10 0
PB3 14 0
PB4 20 0
PB5 24 0

J1 1 2 250u
J2 4 5 200u
J3 4 6 202u
J4 8 9 250u
J5 11 12 200u
J6 11 13 202u
J7 7 15 196u
J8 16 17 165u
J9 18 19 250u
J10 21 16 146u
J11 22 23 250u

.end
