* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===
* Back-annotated simulation file written by InductEx v.6.0.4 on 26-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 26 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			  a q0 q1
.subckt LSMITLL_SPLITT a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param Lptl=2p
.param BiasCoef=0.7
.param RD=1.36

.param B1=1.6
.param B2=1.67
.param B3=2.5
.param B4=2.5
.param IB1=225u
.param IB2=185u
.param IB3=185u
.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))/2
.param L3=(Phi0/(2*B1*Ic0))/2
.param L4=(Phi0/(2*B2*Ic0))/2
.param L5=(Phi0/(2*B2*Ic0))/2
.param L6=Lptl
.param L7=(Phi0/(2*B2*Ic0))/2
.param L8=Lptl
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 8 pwl(0 0 5p IB2)
IB3 0 11 pwl(0 0 5p IB3)
B1 2 3 jjmit area=B1
B2 5 6 jjmit area=B2
B3 8 9 jjmit area=B3
B4 11 12 jjmit area=B4
L1 a 2 1.515E-12
L2 2 4 2.836E-12
L3 4 5 2.85E-12
L4 5 7 2.68E-12
L5 7 8 2.699E-12
L6 8 10 2.364E-12
L7 7 11 2.704E-12
L8 11 13 2.369E-12
LP1 3 0 4.521E-13
LP2 6 0 5.395E-13
LP3 9 0 5.061E-13
LP4 12 0 5.078E-13
RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 5 105 RB2
LRB2 105 0 LRB2
RB3 8 108 RB3
LRB3 108 0 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
RD1 13 q0 RD
RD2 10 q1 RD
.ends

* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 22
b1    1  2  jjmitll100 area=2.25
b2    3  4  jjmitll100 area=2.25
b3    5  6  jjmitll100 area=2.5
ib1   0  2  pwl(0 0 5p 275ua)
ib2   0  5  pwl(0 0 5p 175ua)
l1    8  7  1p
l2    7  0  3.9p
l3    7  1  0.6p
l4    2  3  1.1p
l5    3  5  4.5p
l6    5  11 2p
lp2   4  0  0.2p
lp3   6  0  0.2p
lrb1  9  2  1p
lrb2  10 4  1p
lrb3  12 6  1p
rb1   1  9  4.31
rb2   3  10 4.31
rb3   5  12 3.88
b01   23 27 jjmitll100 area=2
b02   24 26 jjmitll100 area=1.62
ib01  0  30 pwl(0      0 5p 0.00023)
ib02  0  31 pwl(0      0 5p 8.2e-005)
l01   11 23 2.5e-012
l02   23 24 3.3e-012
l03   24 25 3.5e-013
lp01  0  27 5e-014
lp02  0  26 1.2e-013
lpr01 23 30 2e-013
lpr02 24 31 1.3e-012
lrb01 27 28 1e-012
lrb02 26 29 1e-012
rb01  28 23 4.85
rb02  29 24 6.3
rins  25 22 1.36
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
tload 2 0 5 0 lossless z0=5 td=10p
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
tload 2 0 5 0 lossless z0=5 td=50p
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  2
b1    1  9  jjmitll100     area=1
b2    4  8  jjmitll100     area=1
b3    5  7  jjmitll100     area=1
ib1   0  10 pwl(0      0 5p 145u)
l1    2  1  0.2p
l2    1  3  4.3p
l3    3  4  4.6p
l4    4  5  6.0p
l5    5  6  1.3p
lp1   0  9  0.34p
lp2   0  8  0.06p
lp3   0  7  0.03p
lpr1  3  10 0.2p
lrb1  9  11 0.5p
lrb2  8  12 1p
lrb3  7  13 1p
rb1   11 1  15.4
rb2   12 4  11.3
rb3   13 5  11.3
rsink 6  0  2
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160ohm, rn=16ohm, icrit=0.1ma)
.ENDS SINKCELL
* ===== MAIN =====
I_a 0 1 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa SOURCECELL 1 2
XLOADINa LOADINCELL 2 3
XLOADOUTq0 LOADOUTCELL 4 5
XSINKOUTq0 SINKCELL 5
XLOADOUTq1 LOADOUTCELL 6 7
XSINKOUTq1 SINKCELL 7
XDUT lsmitll_splitt 3 4 6
.tran 0.025p 1000p 0
.print i(L1.XDUT) p(B1.XDUT) i(L8.XDUT) p(B4.XDUT) i(L6.XDUT) p(B3.XDUT)
.end
