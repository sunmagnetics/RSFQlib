* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 17 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_OR2T_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 [L1]			
L2 1 4 6.7019p [L2]	
L3 4 7 6.2519p [L3]	
L4 9 10 0.7723p [L4]	
L5 b 11 [L5]
L6 11 14 6.7019p [L6]
L7 14 17 6.2519p [L7]
L8 19 10 0.7723p [L8]
L9 10 21 4.6089p [L9]
L10 22 25 7.7141p [L10]
L11 clk 26 [L11]
L12 26 28 2.7407p [L12]
L13 28 30 3.4070p [L13]
L14 30 32 4.5212p [L14]
L15 25 34 4.5560p [L15]
L16 34 q [L16]

LB1 1 3 [LB1]
LB2 4 6 [LB2]
LB3 11 13 [LB3]
LB4 14 16 [LB4]	
LB5 10 20 [LB5]
LB6 22 24 [LB6]	
LB7 28 29 [LB7]
LB8 34 36 [LB8]	

LP1 2 0 [LP1]
LP2 5 0 [LP2]		
LP3 8 0 [LP3]	
LP5 12 0 [LP5]	
LP6 15 0 [LP6]
LP7 18 0 [LP7]
LP10 23 0 [LP10]	
LP11 27 0 [LP11]	
LP12 31 0 [LP12]	
LP14 33 0 [LP14]
LP15 35 0 [LP15]
	
* Ports
P1 a 0
P2 b 0
P3 clk 0
P4 q 0

PB1 3 0
PB2 6 0
PB3 13 0
PB4 16 0
PB5 20 0
PB6 24 0
PB7 29 0
PB8 36 0

J1 1 2 160u
J2 4 5 128u
J3 7 8 165u
J4 7 9 125u
J5 11 12 160u
J6 14 15 128u
J7 17 18 165u
J8 17 19 125u
J9 21 22 167u
J10 22 23 195u
J11 26 27 160u
J12 30 31 159u
J13 32 25 144u
J14 25 33 209u
J15 34 35 250u

.end