* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 22 June 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_ptlrx_v2p1_base.cir
.endc

* Inductors
L1 a 1 [L1]
L2 1 4 6.37p [L2]
L3 4 7 5.17p [L3]
L4 7 q 2.07p [L4]

LB1 1 3 [LB1]
LB2 4 6 [LB2]
LB3 7 9 [LB3]
LP1 2 0 [LP1]
LP2 5 0 [LP2]
LP3 8 0 [LP3]
* Ports
P1 a 0
P2 q 0
PB1 3 0
PB2 6 0
PB3 9 0
J1 1 2 162u
J2 4 5 200u
J3 7 8 250u
.end