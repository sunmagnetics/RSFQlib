* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 22 June 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_ptltx_v2p1_base.cir
.endc

* Inductors
L1 a 1 2.07p [L1]
L2 1 4 4.14p [L2]
L3 4 7 [L3]
LP1 2 0 [LP1]
LP2 5 0 [LP2]
LB1 1 3 [LB1]
LB2 4 6 [LB2]
* Ports
P1 a 0
P2 7 0
PB1 3 0
PB2 6 0
J1 1 2 250u
J2 4 5 250u
.end