* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 27 April 2021
* Last modification by: L. Schindler

.control
	back-annotate LSmitll_SFQDC_v2p1_base.cir
.endc

* Inductors
L1 1 2 1.522p [L1]
L3 2 5 0.827p [L3]
L4 5 6 1.12884p [L4]
L5 5 7 1.11098p [L5]
L5b 10 12 3.216p [L5b]
L6 8 12 5.94p [L6]
L10 12 17 0.215p [L10]
L19 18 20 0.954p [L19]
L13 20 22 3.699p [L13]
L18 22 24 2.010p [L18]
L17 24 26 1.510p [L17]
LR1 12 13 0.91p [LR1]
LB1 2 3 [LB1]
LB2 8 9 [LB2]
LB3 18 19 [LB3]
LB4 22 23 [LB4]
LP1 4 0 [LP1]
LP4 11 0 [LP4]
LP5 15 0 [LP5]
LP7 21 0 [LP7]
LP8 25 0 [LP8]
* Ports
P1 1 0
P2 3 0
P3 9 0
P4 13 0
P5 19 0
P6 23 0
P7 26 0
J1 2 4 325u
J2 7 10 200u
J3 6 8 150u
J4 10 11 300u
J5 8 15 175u
J6 17 18 150u
J7 20 21 150u
J8 24 25 200u
.end