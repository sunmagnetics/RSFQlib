* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 15 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_PTLTX_v3p0_base.cir
.endc

* Inductors
L1 a 1 2.0678p [L1]
L2 1 4 4.1357p [L2]
L3 4 7 [L3]

LP1 2 0 [LP1]
LP2 5 0 [LP2]

LB1 1 3 [LB1]
LB2 4 6 [LB2]

* Ports
P1 a 0
P2 7 0

PB1 3 0
PB2 6 0

J1 1 2 250u
J2 4 5 250u

.end