* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 6 September 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_XORT_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 [L1]			
L2 1 3 2.7271p [L2]	
L3 3 5 3.7490p [L3]	
L4 5 7 3.4856p [L4]	
L5 9 10 11.3746p [L5]
L6 b 11 [L6]
L7 11 13 2.7271p [L7]
L8 13 15 3.7490p [L8]
L9 15 17 3.4856p [L9]
L10 10 19 11.3746p [L10]
L11 10 21 1.0849p [L11]
L12 clk 24 [L12]
L13 24 26 1.8920p [L13]
L14 26 28 2.9216p [L14]
L15 28 30 4.4126p [L15]
L16 22 31 5.1623p [L16]
L17 31 q [L17]

LB1 4 3 [LB1]
LB2 14 13 [LB2]
LB3 20 10 [LB3]
LB4 27 26 [LB4]	
LB5 33 31 [LB5]

LP1 2 0 [LP1]
LP2 6 0 [LP2]		
LP3 8 0 [LP3]	
LP5 12 0 [LP5]	
LP6 16 0 [LP6]
LP7 18 0 [LP7]
LP10 23 0 [LP10]	
LP11 25 0 [LP11]	
LP12 29 0 [LP12]
LP14 32 0 [LP14]
	
* Ports
P1 a 0
P2 b 0
P3 clk 0
P4 q 0

PB1 4 0
PB2 14 0
PB3 20 0
PB4 27 0
PB5 33 0

J1 1 2 160u
J2 5 6 125u
J3 7 8 245u
J4 7 9 222u
J5 11 12 160u
J6 15 16 125u
J7 17 18 245u
J8 17 19 222u
J9 21 22 156u
J10 22 23 152u
J11 24 25 160u
J12 28 29 216u
J13 30 22 147u
J14 31 32 250u

.end