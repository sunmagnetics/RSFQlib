* Author: L. Schindler
* Version: 1.1.40
* Last modification date: 15 April 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

* Ports 			IN OUT	
.subckt LSmitll_PTLRX a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
B0 3 8 14 jjmit area=1
B1 4 10 15 jjmit area=1
B2 5 12 16 jjmit area=1
I0 0 6 pwl(0 0 5p 155u)
L0 6 7 0.2p
L1 a 3 0.2p
L2 3 7 4.3p
L3 7 4 4.6p
L4 4 5 5p
L5 5 q 2.3p
L6 8 0 0.34p
L7 9 0 0.5p
L8 10 0 0.06p
L9 11 0 1p
L10 12 0 0.03p
L11 13 0 1p
R0 3 9 6.859904418
R1 4 11 6.859904418
R2 5 13 6.859904418
.ends LSmitll_PTLRX