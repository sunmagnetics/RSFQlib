* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 7 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_OR2_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 1.6049e-12 [L1]
L2 1 4 4.4173e-12 [L2]
L3 6 7 0.7163E-12 [L3]
L4 b 8 1.6049e-12 [L4]
L5 8 11 4.4173e-12 [L5]
L6 13 7 0.7163E-12 [L6]
L7 7 15 3.2947e-12 [L7]
L8 16 19 8.7190e-12 [L8]
L9 clk 21 2.1422e-12 [L9]
L10 21 24 3.7843e-12 [L10]
L11 19 25 3.9628e-12 [L11]
L12 25 q 1.6906e-12 [L12]

LB1 1 3 
LB2 8 10 
LB3 7 14 
LB4 16 18 
LB5 23 21 
LB6 25 27 

LP1 2 0 [LP1]
LP2 5 0 [LP2]
LP4 9 0 [LP4]
LP5 12 0 [LP5]
LP8 17 0 [LP8]
LP9 20 0 [LP9]
LP10 22 0 [LP10]
LP12 26 0 [LP12]

* Ports
P1 a 0
P2 b 0
P3 clk 0
P4 q 0

J1 1 2 250u
J2 4 5 167u
J3 4 6 148u
J4 8 9 250u
J5 11 12 167u
J6 11 13 148u
J7 15 16 227u
J8 16 17 236u
J9 19 20 176u
J10 21 22 250u
J11 24 19 144u
J12 25 26 250u

PB1 3 0
PB2 10 0
PB3 14 0
PB4 18 0
PB5 23 0
PB6 27 0
.ends