* Back-annotated simulation file written by InductEx v.6.0.4 on 16-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 3 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports  a b clk q
.subckt LSMITLL_XNOR a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=2.66
.param B3=2.34
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=2.31
.param B8=3.15
.param B9=2.5
.param B10=2.58
.param B11=1.44
.param B12=2.60
.param B13=2.71
.param B14=1.63
.param B15=0.95
.param B16=1.44
.param B17=1.40
.param B18=2.5

.param IB1=175E-6
.param IB2=153E-6
.param IB3=IB1
.param IB4=IB2
.param IB5=175E-6
.param IB6=260E-6
.param IB7=56E-6
.param IB8=248E-6
.param IB9=51E-6
.param IB10=175E-6

.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=1p
.param L4=Phi0/(B2*Ic0)
.param L5=L1
.param L6=L2
.param L7=L3
.param L8=L4
.param L9=1p
.param L10=Lptl
.param L11=Phi0/(2*B9*Ic0)
.param L12=1p
.param L13=1p
.param L14=Phi0/(2*B10*Ic0)
.param L15=Phi0/(4*B12*Ic0)
.param L16=Phi0/(4*B12*Ic0)
.param L17=Phi0/(B13*Ic0)
.param L18=1p
.param L20=1p
.param L21=0.5p
.param L22=Phi0/(B16*Ic0)
.param L23=Phi0/(4*B16*Ic0)
.param L24=Phi0/(2*B17*Ic0)
.param L25=Lptl

.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param RB16=B0Rs/B16
.param RB17=B0Rs/B17
.param RB18=B0Rs/B18
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet
.param LRB16=(RB16/Rsheet)*Lsheet
.param LRB17=(RB17/Rsheet)*Lsheet
.param LRB18=(RB18/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 3 4 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 10 11 jjmit area=B5
B6 12 13 jjmit area=B6
B7 14 15 jjmit area=B7
B8 15 16 jjmit area=B8
B9 17 18 jjmit area=B9
B10 19 20 jjmit area=B10
B11 22 15 jjmit area=B11
B12 23 24 jjmit area=B12
B13 26 27 jjmit area=B13
B14 29 34 jjmit area=B14
B15 34 31 jjmit area=B15
B16 28 33 jjmit area=B16
B17 35 36 jjmit area=B17
B18 37 38 jjmit area=B18

LP1 2 0 5.29E-13
LP2 4 0 4.956E-13
LP4 9 0 4.424E-13
LP5 11 0 5.101E-13
LP8 16 0 5.051E-13
LP9 18 0 5.321E-13
LP10 20 0 5.07E-13
LP12 24 0 5.287E-13
LP13 27 0 5.393E-13
LP17 36 0 5.753E-13
LP18 38 0 5.361E-13

IB1 0 1 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 8 pwl(0 0 5p IB3)
IB4 0 13 pwl(0 0 5p IB4)
IB5 0 17 pwl(0 0 5p IB5)
IB6 0 19 pwl(0 0 5p IB6)
IB7 0 25 pwl(0 0 5p IB7)
IB8 0 34 pwl(0 0 5p IB8)
IB9 0 35 pwl(0 0 5p IB9)
IB10 0 37 pwl(0 0 5p IB10)

L1 a 1 2.058E-12
L2 1 3 2.395E-12
L3 3 5 1.108E-12
L4 6 7 4.1E-12
L5 b 8 2.104E-12
L6 8 10 2.374E-12
L7 10 12 9.887E-13
L8 13 7 4.048E-12
L9 7 14 1.15E-12
L10 clk 17 2.041E-12
L11 17 19 3.442E-12
L12 19 21 8.703E-13
L13 21 22 1.117E-12
L14 21 23 2.107E-12
L15 23 25 1.641E-12
L16 25 26 1.335E-12
L17 26 28 5.203E-12
L18 15 29 1.494E-12
L20 31 32 2.081E-12
L21 33 32 9.13E-13
L22 34 28 6.448E-12
L23 32 35 1.012E-12
L24 35 37 3.546E-12
L25 37 q 2.034E-12

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 3 103 RB2
LRB2 103 0 LRB2
RB3 5 105 RB3
LRB3 105 6 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 10 110 RB5
LRB5 110 0 LRB5
RB6 12 112 RB6
LRB6 112 13 LRB6
RB7 14 114 RB7
LRB7 114 15 LRB7
RB8 15 115 RB8
LRB8 115 0 LRB8
RB9 17 117 RB9
LRB9 117 0 LRB9
RB10 19 119 RB10
LRB10 119 0 LRB10
RB11 22 122 RB11
LRB11 122 15 LRB11
RB12 23 123 RB12
LRB12 123 0 LRB12
RB13 26 126 RB13
LRB13 126 0 LRB13
RB14 29 129 RB14
LRB14 129 34 LRB14
RB15 34 130 RB15
LRB15 130 31 LRB15
RB16 28 128 RB16
LRB16 128 33 LRB16
RB17 35 135 RB17
LRB17 135 0 LRB17
RB18 37 137 RB18
LRB18 137 0 LRB18
.ends
