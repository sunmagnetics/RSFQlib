* Author: L. Schindler
* Version: 1.1.40
* Last modification date: 30 January 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

* Ports 			IN IN CLK OUT	
.subckt LSmitll_OR2T a b clk q
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01=1.9518 
.param B01rx2=1.1720 
.param B01rx3=0.8056 
.param B01tx1=1.9004 
.param B02=1.3074 
.param B02rx3=0.7521 
.param B03rx3=0.6339 
.param B05=1.7221 
.param B08=1.3953 
.param B09=1.6170 
.param B10=2.2048 
.param IB01=0.0003277005 
.param IB01rx2=0.0001412752 
.param IB01rx3=9.8325e-05 
.param IB01tx1=0.0001765029 
.param IB02=8.1358e-05 
.param IB04=8.0964e-05 
.param L01=2.6809e-12 
.param L01rx2=2.0307e-12 
.param L01rx3=1.4136e-12 
.param L01tx1=4.2904e-12 
.param L02=1.3486e-12 
.param L02rx2=2.0822e-12 
.param L02rx3=3.3652e-12 
.param L02tx1=2.7779e-12 
.param L03rx3=4.0267e-12 
.param L05=3.7250e-13 
.param L06=1.8890e-12 
.param L07=2.1922e-13 
.param L08=5.4916e-12 
.param L09=1.5727e-12 
.param L13=2.0776e-12 
.param L14=8.8496e-13 
.param LRB01=(RB01/Rsheet)*Lsheet
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01rx2=(RB01rx2/Rsheet)*Lsheet
.param LRB01rx3=(RB01rx3/Rsheet)*Lsheet
.param LRB01tx1=(RB01tx1/Rsheet)*Lsheet
.param LRB02=(RB02/Rsheet)*Lsheet
.param LRB02rx3=(RB02rx3/Rsheet)*Lsheet
.param LRB03=(RB03/Rsheet)*Lsheet
.param LRB03rx3=(RB03rx3/Rsheet)*Lsheet
.param LRB04=(RB04/Rsheet)*Lsheet
.param LRB05=(RB05/Rsheet)*Lsheet
.param LRB08=(RB08/Rsheet)*Lsheet
.param LRB09=(RB09/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param RB01=B0Rs/B01
.param RB01rx1=B0Rs/B01rx2
.param RB01rx2=B0Rs/B01rx2
.param RB01rx3=B0Rs/B01rx3
.param RB01tx1=B0Rs/B01tx1
.param RB02=B0Rs/B02
.param RB02rx3=B0Rs/B02rx3
.param RB03=B0Rs/B01
.param RB03rx3=B0Rs/B03rx3
.param RB04=B0Rs/B02
.param RB05=B0Rs/B05
.param RB08=B0Rs/B08
.param RB09=B0Rs/B09
.param RB10=B0Rs/B10
B01 7 36 62 jjmit area=B01
B01rx1 9 34 61 jjmit area=B01rx2
B01rx2 19 54 70 jjmit area=B01rx2
B01rx3 6 23 59 jjmit area=B01rx3
B01tx1 16 50 68 jjmit area=B01tx1
B02 7 8 60 jjmit area=B02
B02rx3 5 20 58 jjmit area=B02rx3
B03 17 56 71 jjmit area=B01
B03rx3 5 13 63 jjmit area=B03rx3
B04 17 18 69 jjmit area=B02
B05 11 44 65 jjmit area=B05
B08 14 46 66 jjmit area=B08
B09 15 48 67 jjmit area=B09
B10 10 11 64 jjmit area=B10
IB01 0 28 pwl(0 0 5p IB01)
IB01rx1 0 26 pwl(0 0 5p IB01rx2)
IB01rx2 0 42 pwl(0 0 5p IB01rx2)
IB01rx3 0 25 pwl(0 0 5p IB01rx3)
IB01tx1 0 32 pwl(0 0 5p IB01tx1)
IB02 0 29 pwl(0 0 5p IB02)
IB04 0 31 pwl(0 0 5p IB04)
L01 27 7 L01
L01rx1 a 9 L01rx2
L01rx2 b 19 L01rx2
L01rx3 clk 6 L01rx3
L01tx1 15 16 L01tx1
L02 8 12 L02
L02rx1 9 27 L02rx2
L02rx2 19 52 L02rx2
L02rx3 6 22 L02rx3
L02tx1 16 43 L02tx1
L03 52 17 L01
L03rx3 22 5 L03rx3
L04 12 18 L02
L05 12 38 L05
L06 38 10 L06
L07 11 39 L07
L08 39 13 L08
L09 13 14 L09
L13 14 40 L13
L14 40 15 L14
LP01 36 0 0.2p
LP01rx1 34 0 3.4e-13
LP01rx2 54 0 3.4e-13
LP01rx3 23 0 3.4e-13
LP01tx1 50 0 5e-14
LP02rx3 20 0 3.4e-13
LP03 56 0 2e-13
LP05 44 0 0.2p
LP08 46 0 1.17e-13
LP09 48 0 1.51e-13
LPIB01 28 38 0.2p
LPIB02 29 39 0.2p
LPIB04 31 40 0.2p
LPR01rx1 26 27 0.2p
LPR01rx2 42 52 0.2p
LPR01rx3 22 25 2e-13
LPR01tx1 32 16 0.2p
LRB01 37 0 LRB01
LRB01rx1 35 0 LRB01rx1
LRB01rx2 55 0 LRB01rx2
LRB01rx3 24 0 LRB01rx3
LRB01tx1 51 0 LRB01tx1
LRB02 33 8 LRB02
LRB02rx3 21 0 LRB02rx3
LRB03 57 0 LRB03
LRB03rx3 30 13 LRB03rx3
LRB04 53 18 LRB04
LRB05 45 0 LRB05
LRB08 47 0 LRB08
LRB09 49 0 LRB09
LRB10 41 11 LRB10
RB01 7 37 RB01
RB01rx1 9 35 RB01rx1
RB01rx2 19 55 RB01rx2
RB01rx3 6 24 RB01rx3
RB01tx1 16 51 RB01tx1
RB02 7 33 RB02
RB02rx3 5 21 RB02rx3
RB03 17 57 RB03
RB03rx3 5 30 RB03rx3
RB04 17 53 RB04
RB05 11 45 RB05
RB08 14 47 RB08
RB09 15 49 RB09
RB10 10 41 RB10
RINStx1 43 q 1.36
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.ends LSmitll_OR2T
