* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/09/01.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 30 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	b	clk	q	
.subckt THmitll_NDROT a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=1.6
.param B2=1.45
.param B3=2.15
.param B4=1.73
.param B5=2.54
.param B6=1.6
.param B7=1.45
.param B8=2.15
.param B9=1.73
.param B10=2.54
.param B11=0.74
.param B12=1.57
.param B13=1.6
.param B14=1.6 
.param B15=1.08
.param B16=2.5

.param IB1=268u
.param IB2=129u
.param IB3=225u
.param IB4=268u
.param IB5=129u
.param IB6=115u
.param IB7=254u
.param IB8=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param LB8=LB

.param L1=Lptl
.param L2=2.3873p
.param L3=2.7660p
.param L4=4.1774p
.param L5=3.2486p
.param L6=3.7241p
.param L7=Lptl
.param L8=2.3873p
.param L9=2.7660p
.param L10=4.1774p
.param L11=3.2486p
.param L12=3.7241p
.param L13=0.8049p
.param L14=0.8860p
.param L15=Lptl
.param L16=2.6122p
.param L17=2.6435p
.param L18=3.5452p
.param L19=4.6837p
.param L20=Lptl

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP8=LP
.param LP10=LP
.param LP12=LP
.param LP13=LP
.param LP14=LP
.param LP16=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param RB16=B0Rs/B16

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet+LP
.param LRB13=(RB13/Rsheet)*Lsheet+LP
.param LRB14=(RB14/Rsheet)*Lsheet+LP
.param LRB15=(RB15/Rsheet)*Lsheet
.param LRB16=(RB16/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 10 11 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 15 16 jjmit  area=B6 
B7 19 20 jjmit  area=B7 
B8 21 22 jjmit  area=B8
B9 24 25 jjmit  area=B9 
B10 25 26 jjmit  area=B10 
B11 14 27 jjmit  area=B11 
B12 30 31 jjmit  area=B12 
B13 32 33 jjmit  area=B13 
B14 36 37 jjmit  area=B14 
B15 38 30 jjmit  area=B15 
B16 39 40 jjmit  area=B16 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)
IB6 0 29 pwl(0 0 5p IB6)
IB7 0 35 pwl(0 0 5p IB7)
IB8 0 41 pwl(0 0 5p IB8)

LB1 4 3 8.139E-013 
LB2 9 7 6.905E-013 
LB3 13 11 2.05E-012 
LB4 18 17 7.93E-013 
LB5 23 21 6.92E-013 
LB6 29 28 2.339E-012 
LB7 35 34 2.399E-012 
LB8 41 39 1.726E-012 

L1 a 1 1.001E-012 
L2 1 3 2.395E-012 
L3 3 5 2.766E-012 
L4 5 7 4.17E-012 
L5 7 10 3.25E-012 
L6 11 14 3.695E-012
L7 b 15 1.003E-012 
L8 15 17 2.401E-012 
L9 17 19 2.779E-012 
L10 19 21 4.183E-012 
L11 21 24 3.255E-012 
L12 25 14 3.713E-012 
L13 27 28 8.093E-013 
L14 28 30 8.804E-013 
L15 clk 32 1.351E-012 
L16 32 34 2.624E-012 
L17 34 36 2.63E-012 
L18 36 38 3.565E-012 
L19 30 39 4.674E-012 
L20 39 42 6.06E-013 

RD 42 q RD  

LP1 2 0 3.626E-013 
LP2 6 0 4.608E-013 
LP3 8 0 3.732E-013 
LP5 12 0 4.072E-013 
LP6 16 0 3.63E-013 
LP7 20 0 4.592E-013 
LP8 22 0 3.742E-013 
LP10 26 0 3.912E-013 
LP12 31 0 4.701E-013 
LP13 33 0 3.832E-013 
LP14 37 0 4.271E-013 
LP16 40 0 3.764E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 10 110 RB4  
LRB4 110 11 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 15 115 RB6  
LRB6 115 0 LRB6 
RB7 19 119 RB7  
LRB7 119 0 LRB7 
RB8 21 121 RB8  
LRB8 121 0 LRB8 
RB9 24 124 RB9  
LRB9 124 25 LRB9 
RB10 25 125 RB10  
LRB10 125 0 LRB10 
RB11 14 127 RB11  
LRB11 127 27 LRB11 
RB12 30 130 RB12  
LRB12 130 0 LRB12 
RB13 32 132 RB13  
LRB13 132 0 LRB13 
RB14 36 136 RB14  
LRB14 136 0 LRB14 
RB15 38 138 RB15  
LRB15 138 30 LRB15 
RB16 39 139 RB16  
LRB16 139 0 LRB16 

.ends
