* Author: L. Schindler
* Version: 2.1
* Last modification date: 7 January 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports  a b clk q
.subckt LSMITLL_AND2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC/1.4
.param B3=IC
.param B4=IC/1.4
.param B5=IC
.param B6=IC/1.4
.param B7=B1
.param B8=B2
.param B9=B3
.param B10=B4
.param B11=B5
.param B12=B6
.param B13=IC
.param B14=IC
.param B15=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=BiasCoef*Ic0*B3
.param IB3=IB1
.param IB4=IB2
.param IB5=BiasCoef*Ic0*B13
.param IB6=BiasCoef*Ic0*B14
.param IB7=BiasCoef*Ic0*B15

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB

.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(B3*Ic0)
.param L4=1p
.param L5=Phi0/(2*B5*Ic0)
.param L6=L1
.param L7=L2
.param L8=L3
.param L9=L4
.param L10=L5
.param L11=Phi0/(4*IC*Ic0)
.param L12=Phi0/(2*B13*Ic0)
.param L13=1p
.param L14=1p
.param L15=Phi0/(4*IC*Ic0)

.param LP1=LP
.param LP3=LP
.param LP5=LP
.param LP7=LP
.param LP9=LP
.param LP11=LP
.param LP13=LP
.param LP14=LP
.param LP15=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet
.param LRB15=(RB15/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 8 11 jjmit area=B5
B6 12 13 jjmit area=B6
B7 14 15 jjmit area=B7
B8 17 18 jjmit area=B8
B9 18 19 jjmit area=B9
B10 21 22 jjmit area=B10
B11 21 23 jjmit area=B11
B12 24 13 jjmit area=B12
B13 25 26 jjmit area=B13
B14 31 32 jjmit area=B14
B15 28 29 jjmit area=B15

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 27 pwl(0 0 5p IB5)
IB6 0 33 pwl(0 0 5p IB6)
IB7 0 30 pwl(0 0 5p IB7)

LB1 3 1 LB1
LB2 7 5 LB2
LB3 16 14 LB3
LB4 20 18 LB4
LB5 27 25 LB5
LB6 30 28 LB6
LB7 33 31 LB7

LP1 2 0 LP1
LP3 6 0 LP3
LP5 11 0 LP5
LP7 15 0 LP7
LP9 19 0 LP9
LP11 23 0 LP11
LP13 26 0 LP13
LP14 32 0 LP14
LP15 29 0 LP15

L1 a 1 L1
L2 1 4 L2
L3 5 8 L3
L4 9 10 L4
L5 8 12 L5
L6 b 14 L6
L7 14 17 L7
L8 18 21 L8
L9 22 10 L9
L10 21 24 L10
L11 clk 25 L11
L12 25 31 L12
L13 31 10 L13
L14 13 28 L14
L15 28 q L15

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 5 105 RB3
LRB3 105 0 LRB3
RB4 8 109 RB4
LRB4 109 9 LRB4
RB5 8 108 RB5
LRB5 108 0 LRB5
RB6 12 112 RB6
LRB6 112 13 LRB6
RB7 14 114 RB7
LRB7 114 0 LRB7
RB8 17 117 RB8
LRB8 117 18 LRB8
RB9 18 118 RB9
LRB9 118 0 LRB9
RB10 21 122 RB10
LRB10 122 22 LRB10
RB11 21 121 RB11
LRB11 121 0 LRB11
RB12 24 124 RB12
LRB12 124 13 LRB12
RB13 25 125 RB13
LRB13 125 0 LRB13
RB14 31 131 RB14
LRB14 131 0 LRB14
RB15 28 128 RB15
LRB15 128 0 LRB15
.ends