* Author: L. Schindler
* Version: 2.1
* Last modification date: 13 August 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			 a clk q
.subckt LSMITLL_ALWAYS0T_sync a clk q
.param L1=2p
.param L2=2p
.param L3=2p
L1 a 1 L1
L2 clk 2 L2
L3 3 q L3
RA 1 0 2
RCLK 2 0 2
RQ 3 0 2
.ends