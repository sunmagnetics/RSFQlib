* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 24 June 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

*$Ports 			  a q0 q1
.subckt LSMITLL_CLKSPLT a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01rx1=1.01
.param B01tx1=1.70 
.param B1=1.70 
.param B2=1.21
.param IB01rx1=0.000135
.param IB01tx1=7.6e-05 
.param IB1=0.000360
.param L01rx1=2.6757035519114777e-13 
.param L02tx1=2.2253212527851025e-12 
.param L1=1.5258529970572481e-12 
.param L2=2.9153847294043574e-12 
.param L3=4.813688043861165e-13 
.param L4=1.2716425006912427e-12 
.param L5=1.2572241510058017e-12 
.param LRB01rx1=(RB01rx1/Rsheet)*Lsheet
.param LRB01tx1=(RB01tx1/Rsheet)*Lsheet
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param RB01rx1=B0Rs/B01rx1
.param RB01tx1=B0Rs/B01tx1
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
B01rx1 6 20 jjmit area=B01rx1
B01tx1 5 16 jjmit area=B01tx1
B01tx2 9 28 jjmit area=B01tx1
B1 7 22  jjmit area=B1
B2 4 14  jjmit area=B2
B3 8 25  jjmit area=B2
IB01rx1 0 12 pwl(0 0 5p IB01rx1)
IB01tx1 0 10 pwl(0 0 5p IB01tx1)
IB01tx2 0 27 pwl(0 0 5p IB01tx1)
IB1 0 13 pwl(0 0 5p IB1)
L01rx1 a 6 L01rx1
L02tx1 5 q0 L02tx1
L02tx2 9 q1 L02tx1
L1 6 7 L1
L2 7 18 L2
L3 18 19 L3
L4 4 19 L4
L5 4 5 L5
L6 19 8 L4
L7 8 9 L5
LP01rx1 20 0 0.34p
LP01tx1 16 0 0.05p
LP01tx2 28 0 0.05p
LP1 22 0 0.2p
LP2 14 0 0.2p
LP3 25 0 0.2p
LPR01rx1 12 6 0.2p
LPR01tx1 10 5 0.2p
LPR01tx2 9 27 0.2p
LPRIB1 13 18 0.2p
LRB01rx1 21 0 LRB01rx1
LRB01tx1 17 0 LRB01tx1
LRB01tx2 29 0 LRB01tx1
LRB1 23 0 LRB1
LRB2 15 0 LRB2
LRB3 26 0 LRB2
RB01rx1 6 21 RB01rx1
RB01tx1 5 17 RB01tx1
RB01tx2 9 29 RB01tx1
RB1 7 23 RB1
RB2 4 15 RB2
RB3 8 26 RB2
.ends