* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/29.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 28 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	b	clk	q
.subckt THmitll_XOR a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=2.0
.param B3=2.02
.param B4=2.5
.param B5=2.0
.param B6=2.02
.param B7=1.96
.param B8=1.65
.param B9=2.5
.param B10=1.46
.param B11=2.5

.param IB1=175u
.param IB2=175u
.param IB3=273u
.param IB4=175u
.param IB5=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param L1=1.5740p
.param L2=3.1407p
.param L3=4.7381p
.param L4=1.5740p
.param L5=3.1407p
.param L6=4.7381p
.param L7=4.7751p
.param L8=1.1983p
.param L9=3.2191p
.param L10=3.7711p
.param L11=1.4703p

.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP8=LP
.param LP9=LP
.param LP11=LP

.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8         
.param RB9=B0Rs/B9         
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 4 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 11 13 jjmit  area=B6 
B7 7 15 jjmit  area=B7 
B8 16 17 jjmit  area=B8 
B9 18 19 jjmit  area=B9 
B10 21 16 jjmit  area=B10 
B11 22 23 jjmit  area=B11 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 24 pwl(0 0 5p IB5)

LB1 3 1 8.314E-013 
LB2 10 8 9.179E-013 
LB3 14 7 3.234E-012 
LB4 20 18 1.047E-012 
LB5 24 22 1.004E-012 

L1 a 1 1.57E-012 
L2 1 4 3.128E-012 
L3 6 7 4.746E-012 
L4 b 8 1.578E-012 
L5 8 11 3.145E-012 
L6 7 13 4.763E-012 
L7 15 16 4.74E-012 
L8 clk 18 1.196E-012 
L9 18 21 3.224E-012 
L10 16 22 3.775E-012 
L11 22 q 1.459E-012 

LP1 2 0 4.215E-013 
LP2 5 0 4.657E-013 
LP4 9 0 3.32E-013 
LP5 12 0 3.87E-013 
LP8 17 0 4.698E-013 
LP9 19 0 3.611E-013 
LP11 23 0 4.394E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 4 106 RB3  
LRB3 106 6 LRB3 
RB4 8 108 RB4  
LRB4 108 0 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 11 113 RB6  
LRB6 113 13 LRB6 
RB7 7 115 RB7  
LRB7 115 15 LRB7 
RB8 16 116 RB8  
LRB8 116 0 LRB8 
RB9 18 118 RB9  
LRB9 118 0 LRB9 
RB10 21 121 RB10  
LRB10 121 16 LRB10 
RB11 22 122 RB11  
LRB11 122 0 LRB11 

.ends
