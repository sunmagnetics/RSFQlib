* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 31 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_NDROT_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 [L1]
L2 1 3 2.3876p [L2]
L3 3 5 2.7660p [L3]
L4 5 7 4.1774p [L4]
L5 7 10 3.2486p [L5]
L6 11 14 3.7241p [L6]
L7 b 15 [L7]
L8 15 17 2.3876p [L8]
L9 17 19 2.7660p [L9]
L10 19 21 4.1774p [L10]
L11 21 24 3.2486p [L11]
L12 25 14 3.7241p [L12]
L13 27 28 0.8049p [L13]
L14 28 30 0.8860p [L14]
L15 clk 32 [L15]
L16 32 34 2.6122p [L16]
L17 34 36 2.6435p [L17]
L18 36 38 3.5452p [L18]
L19 30 39 4.6837p [L19]
L20 39 q [L20]

LP1 2 0 [LP1]
LP2 6 0 [LP2]
LP3 8 0 [LP3]
LP5 12 0 [LP5]
LP6 16 0 [LP6]
LP7 20 0 [LP7]
LP8 22 0 [LP8]
LP10 26 0 [LP10]
LP12 31 0 [LP12]
LP13 33 0 [LP13]
LP14 37 0 [LP14]
LP16 40 0 [LP16]

LB1 4 3 [LB1]
LB2 9 7 [LB2]
LB3 13 11 [LB3]
LB4 18 17 [LB4]
LB5 23 21 [LB5]
LB6 29 28 [LB6]
LB7 35 34 [LB7]
LB8 41 39 [LB8]

* Ports
P1 a 0
P2 b 0
P3 clk 0
P4 q 0

PB1 4 0
PB2 9 0
PB3 13 0
PB4 18 0
PB5 23 0
PB6 29 0
PB7 35 0
PB8 41 0

J1 1 2 160u
J2 5 6 145u
J3 7 8 215u
J4 10 11 173u
J5 11 12 254u
J6 15 16 160u
J7 19 20 145u
J8 21 22 215u
J9 24 25 173u
J10 25 26 254u
J11 14 27 74u
J12 30 31 157u
J13 32 33 160u
J14 36 37 160u
J15 38 30 108u
J16 39 40 250u

.end