* Author: L. Schindler
* Version: 3.0
* Last modification date: 30 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	b	clk	q	
.subckt THmitll_NDROT a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=ICreceive
.param B2=IC/1.25
.param B3=IC 
.param B4=IC/1.4
.param B5=IC
.param B6=B1
.param B7=B2
.param B8=B3
.param B9=B4
.param B10=B5
.param B11=IC/3
.param B12=IC/1.25
.param B13=ICreceive
.param B14=IC/1.25 
.param B15=IC/3
.param B16=ICtrans

.param IB1=BiasCoef*Ic0*(B1+B2)
.param IB2=BiasCoef*Ic0*B3
.param IB3=Ic0*B5
.param IB4=IB1
.param IB5=IB2
.param IB6=BiasCoef*Ic0*B12
.param IB7=BiasCoef*Ic0*(B13+B14)
.param IB8=BiasCoef*Ic0*B16

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param LB8=LB

.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))*(B1/(B1+B2))
.param L3=(Phi0/(2*B2*Ic0))*(B2/(B1+B2))
.param L4=Phi0/(2*B2*Ic0)
.param L5=Phi0/(2*B3*Ic0)
.param L6=Phi0/(2*B5*Ic0)
.param L7=Lptl
.param L8=L2
.param L9=L3
.param L10=L4
.param L11=L5
.param L12=L6
.param L13=1p
.param L14=1p
.param L15=Lptl
.param L16=(Phi0/(2*B13*Ic0))*(B13/(B13+B14))
.param L17=(Phi0/(2*B13*Ic0))*(B14/(B13+B14))
.param L18=Phi0/(2*B14*Ic0)
.param L19=Phi0/(2*B12*Ic0)
.param L20=Lptl

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP8=LP
.param LP10=LP
.param LP12=LP
.param LP13=LP
.param LP14=LP
.param LP16=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param RB16=B0Rs/B16

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet+LP
.param LRB13=(RB13/Rsheet)*Lsheet+LP
.param LRB14=(RB14/Rsheet)*Lsheet+LP
.param LRB15=(RB15/Rsheet)*Lsheet
.param LRB16=(RB16/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 10 11 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 15 16 jjmit  area=B6 
B7 19 20 jjmit  area=B7 
B8 21 22 jjmit  area=B8
B9 24 25 jjmit  area=B9 
B10 25 26 jjmit  area=B10 
B11 14 27 jjmit  area=B11 
B12 30 31 jjmit  area=B12 
B13 32 33 jjmit  area=B13 
B14 36 37 jjmit  area=B14 
B15 38 30 jjmit  area=B15 
B16 39 40 jjmit  area=B16 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)
IB6 0 29 pwl(0 0 5p IB6)
IB7 0 35 pwl(0 0 5p IB7)
IB8 0 41 pwl(0 0 5p IB8)

LB1 4 3 LB1 
LB2 9 7 LB2 
LB3 13 11 LB3 
LB4 18 17 LB4 
LB5 23 21 LB5 
LB6 29 28 LB6 
LB7 35 34 LB7 
LB8 41 39 LB8 

L1 a 1 L1 
L2 1 3 L2 
L3 3 5 L3 
L4 5 7 L4 
L5 7 10 L5 
L6 11 14 L6
L7 b 15 L7 
L8 15 17 L8 
L9 17 19 L9 
L10 19 21 L10 
L11 21 24 L11 
L12 25 14 L12 
L13 27 28 L13 
L14 28 30 L14 
L15 clk 32 L15 
L16 32 34 L16 
L17 34 36 L17 
L18 36 38 L18 
L19 30 39 L19 
L20 39 42 L20 

RD 42 q RD  

LP1 2 0 LP1 
LP2 6 0 LP2 
LP3 8 0 LP3 
LP5 12 0 LP5 
LP6 16 0 LP6 
LP7 20 0 LP7 
LP8 22 0 LP8 
LP10 26 0 LP10 
LP12 31 0 LP12 
LP13 33 0 LP13 
LP14 37 0 LP14 
LP16 40 0 LP16 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 10 110 RB4  
LRB4 110 11 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 15 115 RB6  
LRB6 115 0 LRB6 
RB7 19 119 RB7  
LRB7 119 0 LRB7 
RB8 21 121 RB8  
LRB8 121 0 LRB8 
RB9 24 124 RB9  
LRB9 124 25 LRB9 
RB10 25 125 RB10  
LRB10 125 0 LRB10 
RB11 14 127 RB11  
LRB11 127 27 LRB11 
RB12 30 130 RB12  
LRB12 130 0 LRB12 
RB13 32 132 RB13  
LRB13 132 0 LRB13 
RB14 36 136 RB14  
LRB14 136 0 LRB14 
RB15 38 138 RB15  
LRB15 138 30 LRB15 
RB16 39 139 RB16  
LRB16 139 0 LRB16 

.ends
