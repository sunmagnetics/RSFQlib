* Author: L. Schindler
* Version: 3.0
* Last modification date: 3 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports 	a	b	clk	q
.subckt THmitll_OR2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param B3=IC/1.4
.param B4=B1
.param B5=B2
.param B6=B3
.param B7=IC/1.4
.param B8=IC
.param B9=IC
.param B10=IC
.param B11=IC/1.4
.param B12=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=IB1
.param IB3=Ic0*IC
.param IB4=Ic0*B8
.param IB5=BiasCoef*Ic0*B10
.param IB6=BiasCoef*Ic0*B12

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB

.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=1p
.param L4=L1
.param L5=L2
.param L6=L3
.param L7=Phi0/(2*B2*Ic0)
.param L8=Phi0/(B8*Ic0)
.param L9=Phi0/(4*B10*Ic0)
.param L10=Phi0/(2*B10*Ic0)
.param L11=Phi0/(2*B9*Ic0)
.param L12=Phi0/(4*B12*Ic0)

.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP8=LP
.param LP9=LP
.param LP10=LP
.param LP12=LP

.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10 
.param RB11=B0Rs/B11 
.param RB12=B0Rs/B12 

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 4 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 11 13 jjmit  area=B6 
B7 15 16 jjmit  area=B7 
B8 16 17 jjmit  area=B8 
B9 19 20 jjmit  area=B9 
B10 21 22 jjmit  area=B10 
B11 24 19 jjmit  area=B11 
B12 25 26 jjmit  area=B12 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
IB5 0 23 pwl(0 0 5p IB5)
IB6 0 27 pwl(0 0 5p IB6)

LB1 3 1 LB1 
LB2 10 8 LB2 
LB3 14 7 LB3 
LB4 18 16 LB4 
LB5 23 21 LB5 
LB6 27 25 LB6 

L1 a 1 L1 
L2 1 4 L2 
L3 6 7 L3 
L4 b 8 L4 
L5 8 11 L5 
L6 13 7 L6 
L7 7 15 L7 
L8 16 19 L8 
L9 clk 21 L9 
L10 21 24 L10 
L11 19 25 L11 
L12 25 q L12 

LP1 2 0 LP1 
LP2 5 0 LP2 
LP4 9 0 LP4 
LP5 12 0 LP5 
LP8 17 0 LP8 
LP9 20 0 LP9 
LP10 22 0 LP10 
LP12 26 0 LP12 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 4 106 RB3  
LRB3 106 6 LRB3 
RB4 8 108 RB4  
LRB4 108 0 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 11 113 RB6  
LRB6 113 13 LRB6 
RB7 15 115 RB7  
LRB7 115 16 LRB7 
RB8 16 116 RB8  
LRB8 116 0 LRB8 
RB9 19 119 RB9  
LRB9 119 0 LRB9 
RB10 21 121 RB10  
LRB10 121 0 LRB10 
RB11 24 124 RB11  
LRB11 124 19 LRB11 
RB12 25 125 RB12  
LRB12 125 0 LRB12 

.ends
