* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 10 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_SPLITT_v3p0_optimised.cir
.endc

* Inductors
L1 a 1 [L1] 
L2 1 3 2.1010p [L2]
L3 3 5 3.6142p [L3]
L4 5 7 1.7400p [L4]
L5 8 7 1.8162P [L5]
L6 8 q0 [L6]    
L7 7 12 1.8162p [L7]
L8 12 q1 [L8]
LP1 2 0 [LP1] 
LP2 6 0 [LP2] 
LP3 9 0 [LP3]
LP4 13 0 [LP4]
LB1 4 3 [LB1]
LB2 10 8 [LB2]
LB3 14 12 [LB3]

* Ports
P1 a 0
P2 q0 0
P3 q1 0
PB1 4 0
PB2 10 0
PB3 14 0
J1 1 2		160u
J2 5 6 		136u
J3 8 9		250u
J4 12 13	250u
.end
