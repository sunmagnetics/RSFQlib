* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

*             in out
*$Ports  				a  q
.subckt LSmitll_bufft  a  q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
B1 2 3 jjmit area=2.0
B2 6 7 jjmit area=2.5
B3 11 12 jjmit area=2.5
IB1 0 5 pwl(0 0 5p 160u)
IB2 0 10 pwl(0 0 5p 350u)
L1 a 2 2p
L2 2 6 5.2p   
L3 6 9 2.07p
L4 9 11 2.07p
L5 11 14 2p
RD 14 q 1.36
LP1 3 0 0.2p
LP2 7 0 0.2p
LP3 12 0 0.2p
RB1 2 4 3.43
RB2 6 8 2.744
RB3 11 13 2.744
LRB1 4 0 1.94p
LRB2 8 0 1.55p
LRB3 13 0 1.55p
LB1 2 5 1p
LB2 9 10 1p
.ends