* Author: L. Schindler
* Version: 1.1.40
* Last modification date: 30 January 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

* Ports 			IN OUT	
.subckt LSmitll_JTLT a q
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B01=0.6979 
.param B05=1.7851 
.param B02=0.4432
.param B03=0.4881
.param IB01=8.6452e-05 
.param IB03=5.5312e-05
.param IB02=0.000120082 
.param L01=3.3252e-13 
.param L02=2.4032e-12 
.param L03=1.6773e-12 
.param L04=2.5109e-12 
.param L05=8.6652e-13 
.param L07=2.3256e-12 
.param L08=2.3630e-12 
.param LRB03=(RB03/Rsheet)*Lsheet
.param LRB04=(RB04/Rsheet)*Lsheet
.param LRB01=(RB01/Rsheet)*Lsheet
.param LRB05=(RB05/Rsheet)*Lsheet
.param LRB02=(RB02/Rsheet)*Lsheet
.param RB01=B0Rs/B01
.param RB05=B0Rs/B05
.param RB02=B0Rs/B02
.param RB03=B0Rs/B03
.param RB04=B0Rs/B03
B01 3 14 24 jjmit area=B01
B02 4 16 25 jjmit area=B02
B03 5 18 26 jjmit area=B03
B04 6 20 27 jjmit area=B03
B05 7 22 28 jjmit area=B05
IB01 0 8 pwl(0 0 5p IB01)
IB02 0 9 pwl(0 0 5p IB02)
IB03 0 10 pwl(0 0 5p IB03)
L01 a 3 L01
L02 3 11 L02
L03 11 4 L03
L04 4 5 L04
L05 5 12 L05
L06 12 6 L05
L07 6 7 L07
L08 7 13 L08
LB01 8 11 2e-13
LB02 9 12 2e-13
LB03 10 7 2e-13
LP01 14 0 2e-13
LP02 16 0 2e-13
LP03 18 0 2e-13
LP04 20 0 2e-13
LP05 22 0 2e-13
LRB01 15 0 LRB01
LRB02 17 0 LRB02
LRB03 19 0 LRB03
LRB04 21 0 LRB04
LRB05 23 0 LRB05
RB01 3 15 RB01
RB02 4 17 RB02
RB03 5 19 RB03
RB04 6 21 RB04
RB05 7 23 RB05
RINStx 13 q 1.36
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.ends LSmitll_jtlt