* Back-annotated simulation file written by InductEx v.6.0.4 on 15-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 9 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports a b clk q
.subckt LSmitll_NDRO a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=1.99
.param B3=2.2
.param B4=2.5
.param B5=2.35
.param B6=3.24
.param B7=0.74
.param B8=2.5
.param B9=1.17
.param B10=1.09
.param B11=2.5

.param IB1=175u
.param IB2=271u
.param IB3=175u
.param IB4=175u
.param IB5=136u
.param IB6=175u

.param L1=Phi0/(4*IC*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B3*Ic0)
.param L4=Phi0/(4*IC*Ic0)
.param L5=Phi0/(2*B4*Ic0)
.param L6=Phi0/(2*B6*Ic0)
.param L7=1p
.param L8=1p
.param L9=Phi0/(4*IC*Ic0)
.param L10=Phi0/(2*B8*Ic0)
.param L11=Phi0/(2*B10*Ic0)
.param L12=Phi0/(4*IC*Ic0)

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB

B1 1 2 jjmit area=B1
B2 3 4 jjmit area=B2
B3 4 5 jjmit area=B3
B4 7 8 jjmit area=B4
B5 9 10 jjmit area=B5
B6 10 11 jjmit area=B6
B7 6 12 jjmit area=B7
B8 14 15 jjmit area=B8
B9 14 16 jjmit area=B9
B10 17 18 jjmit area=B10
B11 19 20 jjmit area=B11

IB1 0 21 pwl(0 0 5p IB1)
IB2 0 22 pwl(0 0 5p IB2)
IB3 0 23 pwl(0 0 5p IB3)
IB4 0 24 pwl(0 0 5p IB4)
IB5 0 25 pwl(0 0 5p IB5)
IB6 0 26 pwl(0 0 5p IB6)

LB1 1 21 LB1
LB2 4 22 LB2
LB3 7 23 LB3
LB4 14 24 LB4
LB5 13 25 LB5
LB6 19 26 LB6

L1 a 1 2.067E-12
L2 1 3 9.786E-13
L3 4 6 2.693E-12
L4 b 7 2.068E-12
L5 7 9 2.319E-12
L6 10 6 3.438E-12
L7 12 13 1.12E-12
L8 13 17 1.028E-12
L9 clk 14 2.106E-12
L10 16 17 3.135E-12
L11 17 19 3.223E-12
L12 19 q 2.071E-12

LP1 2 0 5.174E-13
LP3 5 0 5.135E-13
LP4 8 0 4.756E-13
LP6 11 0 4.841E-13
LP8 15 0 4.705E-13
LP10 18 0 5.961E-13
LP11 20 0 4.832E-13

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 3 103 RB2
LRB2 103 4 LRB2
RB3 4 104 RB3
LRB3 104 0 LRB3
RB4 7 107 RB4
LRB4 107 0 LRB4
RB5 9 109 RB5
LRB5 109 10 LRB5
RB6 10 110 RB6
LRB6 110 0 LRB6
RB7 6 106 RB7
LRB7 106 12 LRB7
RB8 14 114 RB8
LRB8 114 0 LRB8
RB9 14 116 RB9
LRB9 116 16 LRB9
RB10 17 117 RB10
LRB10 117 0 LRB10
RB11 19 119 RB11
LRB11 119 0 LRB11
.ends
