* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/10.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 10 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$Ports 	a	q0	q1
.subckt THmitll_SPLITT a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=1.6
.param B2=1.36
.param B3=2.5
.param B4=2.5

.param IB1=231u
.param IB2=175u
.param IB3=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB

.param L1=Lptl
.param L2=2.1010p
.param L3=3.6142p
.param L4=1.7400p
.param L5=1.8162p
.param L6=Lptl
.param L7=1.8162p
.param L8=Lptl

.param RD1=RD
.param RD2=RD

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP4=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 8 9 jjmit  area=B3 
B4 12 13 jjmit  area=B4 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 10 pwl(0 0 5p IB2)
IB3 0 14 pwl(0 0 5p IB3)

LB1 4 3 4.087E-013 
LB2 10 8 1.617E-012 
LB3 14 12 2.099E-012 

L1 a 1 1.432E-012 
L2 1 3 2.097E-012 
L3 3 5 3.589E-012 
L4 5 7 1.755E-012 
L5 8 7 1.82E-012 
L6 8 11 7.505E-013 
L7 7 12 1.805E-012 
L8 12 15 1.137E-012 

RD1 11 q0 RD1  
RD2 15 q1 RD2  

LP1 2 0 3.952E-013 
LP2 6 0 4.754E-013 
LP3 9 0 3.421E-013 
LP4 13 0 3.856E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 8 108 RB3  
LRB3 108 0 LRB3 
RB4 12 112 RB4  
LRB4 112 0 LRB4 

.ends

