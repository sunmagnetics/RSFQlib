* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/25.
* Author: T. Hall
* Version: 3.0
* Last modification date: 24 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports 	a	clk	q
.subckt THmitll_NOT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=0.78
.param B3=0.85
.param B4=2.69
.param B5=2.5
.param B6=1.42
.param B7=1.01
.param B8=2.5

.param IB1=175u
.param IB2=131u
.param IB3=175u
.param IB4=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB

.param L1=0.8555p
.param L2=2.7537p
.param L3=0.7553p
.param L4=7.3609p
.param L5=0.8585p
.param L6=3.0349p
.param L7=0.9373p
.param L8=4.2782p
.param L9=0.9209p

.param LP1=LP
.param LP5=LP
.param LP7=LP
.param LP8=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 9 10 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 10 14 jjmit  area=B6 
B7 8 15 jjmit  area=B7 
B8 16 17 jjmit  area=B8 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)

LB1 3 1 1.246E-012 
LB2 6 5 1.707E-012 
LB3 13 11 8.002E-013 
LB4 18 16 8.582E-013 

L1 a 1 8.521E-013 
L2 1 4 2.756E-012 
L3 5 7 7.55E-013 
L4 5 9 7.358E-012 
L5 clk 11 8.595E-013 
L6 11 10 3.051E-012 
L7 8 14 9.435E-013 
L8 8 16 4.287E-012 
L9 16 q 9.3E-013 

LP1 2 0 3.288E-013 
LP5 12 0 3.499E-013 
LP7 15 0 4.831E-013 
LP8 17 0 3.407E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 5 LRB2 
RB3 7 107 RB3  
LRB3 107 8 LRB3 
RB4 9 109 RB4  
LRB4 109 10 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 10 110 RB6  
LRB6 110 14 LRB6 
RB7 8 108 RB7  
LRB7 108 0 LRB7 
RB8 16 116 RB8  
LRB8 116 0 LRB8 

.ends
