* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 2.1
* Last modification date: 18 January 2021
* Last modification by: L. Schindler

* Inductors
L1 1 2 
L2 2 5 2.1p
L3 5 7 1p
L4 8 10 4.12p
L5 11 12 
L6 12 15 2.1p
L7 15 17 1p
L8 18 10 4.12p
L9 10 20 1p
L10 23 24 
L11 24 27 3.11p
L12 27 30 1.07p
L13 31 21 1.01p
L14 30 32 2.45p
L15 32 34 1.83p
L16 34 36 1.12p
L17 36 38 4.32p
L18 21 39 1.6p
L20 42 44 1.06p
L21 43 44 0.55p
L22 38 40 5.40p
L23 44 45 1.18p
L24 45 48 2.78p
L25 48 51 

LB1 2 4
LB2 8 9
LB3 12 14
LB4 18 19
LB5 24 26
LB6 27 29
LB7 34 35
LB8 40 41
LB9 45 47
LB10 48 50

LP1 3 0 
LP2 6 0 
LP4 13 0 
LP5 16 0
LP8 22 0
LP9 25 0 
LP10 28 0
LP12 33 0
LP13 37 0
LP17 46 0
LP18 49 0

* Ports
P1 1 0
P2 11 0
P3 23 0
P4 51 0

PB1 4 0
PB2 9 0
PB3 14 0
PB4 19 0
PB5 26 0
PB6 29 0
PB7 35 0
PB8 41 0
PB9 47 0
PB10 50 0

J1 2 3 200
J2 5 6 274
J3 7 8 223
J4 12 13 200
J5 15 16 274
J6 17 18 223
J7 20 21 240
J8 21 22 329
J9 24 25 200
J10 27 28 242
J11 30 31 136
J12 32 33 240
J13 36 37 228
J14 39 40 175
J15 40 42 107
J16 38 43 154
J17 45 46 164
J18 48 49 250
.end