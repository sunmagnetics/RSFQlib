* Author: L. Schindler
* Version: 3.0
* Last modification date: 30 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports 	a	b	clk	q
.subckt THmitll_NDRO a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC/1.4
.param B3=IC
.param B4=IC
.param B5=IC/1.4
.param B6=IC
.param B7=IC/3
.param B8=IC
.param B9=IC
.param B10=IC/1.4
.param B11=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=Ic0*B3
.param IB3=BiasCoef*Ic0*B4
.param IB4=BiasCoef*Ic0*B8
.param IB5=BiasCoef*Ic0*B9
.param IB6=BiasCoef*Ic0*B11

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB

.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B3*Ic0)
.param L4=Phi0/(4*B4*Ic0)
.param L5=Phi0/(2*B4*Ic0)
.param L6=Phi0/(2*B6*Ic0)
.param L7=2p
.param L8=2p
.param L9=Phi0/(4*B9*Ic0)
.param L10=Phi0/(2*B9*Ic0)
.param L11=Phi0/(2*B8*Ic0)
.param L12=Phi0/(4*B11*Ic0)

.param LP1=LP
.param LP3=LP
.param LP4=LP
.param LP6=LP
.param LP8=LP
.param LP9=LP
.param LP11=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 5 6 jjmit  area=B3 
B4 9 10 jjmit  area=B4 
B5 12 13 jjmit  area=B5 
B6 13 14 jjmit  area=B6 
B7 8 15 jjmit  area=B7 
B8 18 19 jjmit  area=B8 
B9 20 21 jjmit  area=B9 
B10 23 18 jjmit  area=B10 
B11 24 25 jjmit  area=B11 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 11 pwl(0 0 5p IB3)
IB4 0 17 pwl(0 0 5p IB4)
IB5 0 22 pwl(0 0 5p IB5)
IB6 0 26 pwl(0 0 5p IB6)

LB1 3 1 LB1 
LB2 7 5 LB2 
LB3 11 9 LB3 
LB4 17 16 LB4 
LB5 22 20 LB5 
LB6 26 24 LB6 

L1 a 1 L1 
L2 1 4 L2 
L3 5 8 L3 
L4 b 9 L4 
L5 9 12 L5 
L6 13 8 L6 
L7 15 16 L7 
L8 16 18 L8 
L9 clk 20 L9 
L10 20 23 L10 
L11 18 24 L11 
L12 24 q L12 

LP1 2 0 LP1 
LP3 6 0 LP3 
LP4 10 0 LP4 
LP6 14 0 LP6 
LP8 19 0 LP8 
LP9 21 0 LP9 
LP11 25 0 LP11 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 5 LRB2 
RB3 5 105 RB3  
LRB3 105 0 LRB3 
RB4 9 109 RB4  
LRB4 109 0 LRB4 
RB5 12 112 RB5  
LRB5 112 13 LRB5 
RB6 13 113 RB6  
LRB6 113 0 LRB6
RB7 8 108 RB7  
LRB7 108 15 LRB7 
RB8 18 118 RB8  
LRB8 118 0 LRB8 
RB9 20 120 RB9  
LRB9 120 0 LRB9 
RB10 23 123 RB10  
LRB10 123 18 LRB10 
RB11 24 124 RB11  
LRB11 124 0 LRB11 

.ends
