* Back-annotated simulation file written by InductEx v.6.0 on 2021/06/22.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 22 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports a q
.subckt LSmitll_PTLRX a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param LB=2p
.param Lptl=2p
.param IC=2.5
.param BiasCoef=0.7

.param B1=IC/1.54
.param B2=IC/1.25
.param B3=IC
.param IB1=Ic0*B1
.param IB2=BiasCoef*Ic0*B2
.param IB3=BiasCoef*Ic0*B3
.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=Phi0/(2*B2*Ic0)
.param L4=Phi0/(4*IC*Ic0)

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LP1=LP         
.param LP2=LP          
.param LP3=LP  
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3   
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 7 8 jjmit area=B3
IB1 0 3 pwl(0 0 5p IB1)
LB1 1 3 2.777E-012
IB2 0 6 pwl(0 0 5p IB2)
LB2 4 6 2.685E-012
IB3 0 9 pwl(0 0 5p IB3)
LB3 7 9 2.764E-012
L1 a 1 1.346E-012
L2 1 4 6.348E-012
L3 4 7 5.197E-012
L4 7 q 2.058E-012

LP1 2 0 4.795E-013
LP2 5 0 5.431E-013
LP3 8 0 5.339E-013
RB1 1 101 RB1
RB2 4 104 RB2
RB3 7 107 RB3
LRB1 101 0 LRB1
LRB2 104 0 LRB2
LRB3 107 0 LRB3
.ends
