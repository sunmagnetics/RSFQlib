* JSIM deck file generated with TimEx
* === DEVICE-UNDER-TEST ===
* Back-annotated simulation file written by InductEx v.6.0.4 on 28-4-21.
* Author: L. Schindler
* Version: 2.1
* Last modification date: 28 April 2021
* Last modification by: L. Schindler
* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University
* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:
* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.
* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.
*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za
*$ports a b clk q
.subckt LSMITLL_OR2T a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param Lptl=2p
.param LB=2p
.param RD=1.36
.param B1=1.17
.param B2=1.95
.param B3=1.31
.param B4=1.17
.param B5=1.95
.param B6=1.31
.param B7=2.20
.param B8=1.72
.param B9=0.81
.param B10=0.75
.param B11=0.63
.param B12=1.40
.param B13=1.62
.param B14=1.9
.param IB1=141u
.param IB2=141u
.param IB3=328u
.param IB4=81u
.param IB5=98u
.param IB6=81u
.param IB7=177u
.param L1=Lptl
.param L2=2.0822p
.param L3=2.6809p
.param L4=1.3486p
.param L5=Lptl
.param L6=2.0822p
.param L7=2.6809p
.param L8=1.3486p 
.param L10=1.8890p
.param L12=5.4916p
.param L13=Lptl
.param L14=3.3652p
.param L15=4.0267p 
.param L16=0.7p
.param L17=1.5727p
.param L18=2.0776p
.param L19=0.885p
.param L20=4.2904p 
.param L21=Lptl
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param LP1=LP
.param LP2=LP
.param LP4=LP
.param LP5=LP
.param LP8=LP
.param LP9=LP
.param LP10=LP
.param LP12=LP
.param LP13=LP
.param LP14=LP
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11   
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet+LP
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
.param LRB12=(RB12/Rsheet)*Lsheet+LP
.param LRB13=(RB13/Rsheet)*Lsheet+LP
.param LRB14=(RB14/Rsheet)*Lsheet+LP
B1 2 3   jjmit area=B1
B2 6 7   jjmit area=B2
B3 6 8  jjmit area=B3
B4 11 12 jjmit area=B4
B5 15 16 jjmit area=B5
B6 15 43 jjmit area=B6
B7 19 22 jjmit area=B7
B8 22 21 jjmit area=B8
B9 26 27 jjmit area=B9
B10 30 31 jjmit area=B10
B11 32 24 jjmit area=B11
B12 33 34 jjmit area=B12
B13 37 38 jjmit area=B13
B14 39 41 jjmit area=B14
IB1 0 5  pwl(0 0 5p IB1)
IB2 0 14 pwl(0 0 5p IB2)
IB3 0 18 pwl(0 0 5p IB3)
IB4 0 23 pwl(0 0 5p IB4)
IB5 0 29 pwl(0 0 5p IB5)
IB6 0 36 pwl(0 0 5p IB6)
IB7 0 40 pwl(0 0 5p IB7)
L1 a 2 1.593E-12  
L2 2 4 2.116E-12 
L3 4 6 2.655E-12 
L4 8 9 1.349E-12 
L5 b 11 1.596E-12   
L6 11 13 2.104E-12 
L7 13 15 2.655E-12  
L8 43 9 1.348E-12  
L10 9 19 1.883E-12 
L12 22 24 5.465E-12 
L13 clk 26 1.54E-12  
L14 26 28 3.367E-12 
L15 28 30 4.045E-12 
L16 30 32 5.696E-13 
L17 24 33 1.584E-12 
L18 33 35 2.075E-12 
L19 35 37 9.15E-13 
L20 37 39 4.26E-12 
L21 39 42 7.721E-13 
RD 42 q RD
LB1 4 5 2.162E-12
LB2 13 14 2.177E-12
LB3 9 18 2.831E-12
LB4 22 23 3.933E-12
LB5 28 29 1.367E-12
LB6 35 36 2.221E-12
LB7 39 40 2.035E-12
LP1 3 0  4.886E-13
LP2 7 0  4.645E-13
LP4 12 0 4.935E-13
LP5 16 0 4.65E-13
LP8 21 0 5.102E-13
LP9 27 0 5.216E-13
LP10 31 0 5.841E-13
LP12 34 0 4.758E-13
LP13 38 0 5.26E-13
LP14 41 0 4.366E-13
RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 6 106 RB2
LRB2 106 0 LRB2
RB3 6 108 RB3
LRB3 108 8 LRB3
RB4 11 111 RB4
LRB4 111 0 LRB4
RB5 15 115 RB5
LRB5 115 0 LRB5
RB6 15 143 RB6
LRB6 143 43 LRB6
RB7 19 119 RB7
LRB7 119 22 LRB7
RB8 22 122 RB8
LRB8 122 0 LRB8
RB9 26 126 RB9
LRB9 126 0 LRB9
RB10 30 130 RB10
LRB10 130 0 LRB10
RB11 32 132 RB11
LRB11 132 24 LRB11
RB12 33 133 RB12
LRB12 133 0 LRB12
RB13 37 137 RB13
LRB13 137 0 LRB13
RB14 39 139 RB14
LRB14 139 0 LRB14
.ends
* === SOURCE DEFINITION ===
.SUBCKT SOURCECELL  8 22
b1    1  2  jjmitll100 area=2.25
b2    3  4  jjmitll100 area=2.25
b3    5  6  jjmitll100 area=2.5
ib1   0  2  pwl(0 0 5p 275ua)
ib2   0  5  pwl(0 0 5p 175ua)
l1    8  7  1p
l2    7  0  3.9p
l3    7  1  0.6p
l4    2  3  1.1p
l5    3  5  4.5p
l6    5  11 2p
lp2   4  0  0.2p
lp3   6  0  0.2p
lrb1  9  2  1p
lrb2  10 4  1p
lrb3  12 6  1p
rb1   1  9  4.31
rb2   3  10 4.31
rb3   5  12 3.88
b01   23 27 jjmitll100 area=2
b02   24 26 jjmitll100 area=1.62
ib01  0  30 pwl(0      0 5p 0.00023)
ib02  0  31 pwl(0      0 5p 8.2e-005)
l01   11 23 2.5e-012
l02   23 24 3.3e-012
l03   24 25 3.5e-013
lp01  0  27 5e-014
lp02  0  26 1.2e-013
lpr01 23 30 2e-013
lpr02 24 31 1.3e-012
lrb01 27 28 1e-012
lrb02 26 29 1e-012
rb01  28 23 4.85
rb02  29 24 6.3
rins  25 22 1.36
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.ENDS SOURCECELL
* === INPUT LOAD DEFINITION ===
.SUBCKT LOADINCELL  2 5
tload 2 0 5 0 lossless z0=5 td=10p
.ENDS LOADINCELL
* === OUTPUT LOAD DEFINITION ===
.SUBCKT LOADOUTCELL  2 5
tload 2 0 5 0 lossless z0=5 td=50p
.ENDS LOADOUTCELL
* === SINK DEFINITION ===
.SUBCKT SINKCELL  2
b1    1  9  jjmitll100     area=1
b2    4  8  jjmitll100     area=1
b3    5  7  jjmitll100     area=1
ib1   0  10 pwl(0      0 5p 145u)
l1    2  1  0.2p
l2    1  3  4.3p
l3    3  4  4.6p
l4    4  5  6.0p
l5    5  6  1.3p
lp1   0  9  0.34p
lp2   0  8  0.06p
lp3   0  7  0.03p
lpr1  3  10 0.2p
lrb1  9  11 0.5p
lrb2  8  12 1p
lrb3  7  13 1p
rb1   11 1  15.4
rb2   12 4  11.3
rb3   13 5  11.3
rsink 6  0  2
.model jjmitll100 jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160ohm, rn=16ohm, icrit=0.1ma)
.ENDS SINKCELL
* ===== MAIN =====
I_a 0 1 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa SOURCECELL 1 2
XLOADINa LOADINCELL 2 3
I_b 0 4 pwl(0 0 350p 0 353p 600u 356p 0 450p 0 453p 600u 456p 0 480p 0 483p 600u 486p 0 560p 0 563p 600u 566p 0 580p 0 583p 600u 586p 0 660p 0 663p 600u 666p 0 740p 0 743p 600u 746p 0)
XSOURCEINb SOURCECELL 4 5
XLOADINb LOADINCELL 5 6
I_clk 0 7 pulse(0 600u 20p 2p 2p 1p 100p)
XSOURCEINclk SOURCECELL 7 8
XLOADINclk LOADINCELL 8 9
XLOADOUTq LOADOUTCELL 10 11
XSINKOUTq SINKCELL 11
XDUT lsmitll_or2t 3 6 9 10
.tran 0.025p 1000p 0
.print i(L1.XDUT) p(B1.XDUT) i(L5.XDUT) p(B4.XDUT) i(L13.XDUT) p(B9.XDUT) i(L21.XDUT) p(B14.XDUT)
.end
