* Author: L. Schindler
* Version: 3.0
* Last modification date: 3 September 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$ports 	a	b	clk	q
.subckt THmitll_XORT a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=ICreceive
.param B2=IC/1.25
.param B3=IC
.param B4=IC
.param B5=B1
.param B6=B2
.param B7=B3
.param B8=B4
.param B9=IC/1.25
.param B10=IC
.param B11=ICreceive
.param B12=IC/1.25
.param B13=IC/1.4
.param B14=ICtrans

.param IB1=BiasCoef*Ic0*(B1+B2)
.param IB2=IB1
.param IB3=BiasCoef*Ic0*(B3+B7+B9)
.param IB4=BiasCoef*Ic0*(B11+B12)
.param IB5=BiasCoef*Ic0*B14

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP10=LP
.param LP11=LP
.param LP12=LP
.param LP14=LP

.param L1=Lptl
.param L2=(Phi0/(2*B1*Ic0))*(B1/(B1+B2))
.param L3=(Phi0/(2*B1*Ic0))*(B2/(B1+B2))
.param L4=Phi0/(2*B2*Ic0)
.param L5=Phi0/(B3*Ic0)
.param L6=L1
.param L7=L2
.param L8=L3
.param L9=L4
.param L10=L5
.param L11=1.2p
.param L12=Lptl
.param L13=(Phi0/(2*B11*Ic0))*(B11/(B11+B12))
.param L14=(Phi0/(2*B11*Ic0))*(B12/(B11+B12))
.param L15=Phi0/(2*B12*Ic0)
.param L16=Phi0/(2*B10*Ic0)
.param L17=Lptl

.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11   
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
.param LRB12=(RB12/Rsheet)*Lsheet+LP
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 7 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 15 16 jjmit  area=B6 
B7 17 18 jjmit  area=B7 
B8 17 19 jjmit  area=B8 
B9 21 22 jjmit  area=B9 
B10 22 23 jjmit  area=B10 
B11 24 25 jjmit  area=B11 
B12 28 29 jjmit  area=B12 
B13 30 22 jjmit  area=B13 
B14 31 32 jjmit  area=B14 

IB1 0 4 pwl(0 0 5p IB1)
IB2 0 14 pwl(0 0 5p IB2)
IB3 0 20 pwl(0 0 5p IB3)
IB4 0 27 pwl(0 0 5p IB4)
IB5 0 33 pwl(0 0 5p IB5)

LB1 4 3 LB1 
LB2 14 13 LB2 
LB3 20 10 LB3 
LB4 27 26 LB4 
LB5 33 31 LB5 

L1 a 1 L1 
L2 1 3 L2 
L3 3 5 L3 
L4 5 7 L4 
L5 9 10 L5 
L6 b 11 L6 
L7 11 13 L7 
L8 13 15 L8 
L9 15 17 L9 
L10 10 19 L10 
L11 10 21 L11 
L12 clk 24 L12 
L13 24 26 L13 
L14 26 28 L14 
L15 28 30 L15 
L16 22 31 L16 
L17 31 34 L17 

RD 34 q RD  

LP1 2 0 LP1 
LP2 6 0 LP2 
LP3 8 0 LP3 
LP5 12 0 LP5 
LP6 16 0 LP6 
LP7 18 0 LP7 
LP10 23 0 LP10 
LP11 25 0 LP11 
LP12 29 0 LP12 
LP14 32 0 LP14 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 7 109 RB4  
LRB4 109 9 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 15 115 RB6  
LRB6 115 0 LRB6 
RB7 17 117 RB7  
LRB7 117 0 LRB7 
RB8 17 119 RB8  
LRB8 119 19 LRB8 
RB9 21 121 RB9  
LRB9 121 22 LRB9 
RB10 22 122 RB10  
LRB10 122 0 LRB10 
RB11 24 124 RB11  
LRB11 124 0 LRB11 
RB12 28 128 RB12  
LRB12 128 0 LRB12 
RB13 30 130 RB13  
LRB13 130 22 LRB13 
RB14 31 131 RB14  
LRB14 131 0 LRB14 

.ends
