* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/07/25.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 25 July 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports a	q0	q1
.subckt THmitll_SPLIT a q0 q1
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=IC
.param B2=IC
.param B3=IC

.param IB1=BiasCoef*Ic0*B1
.param IB2=BiasCoef*Ic0*B2
.param IB3=IB2

.param LB1=LB
.param LB2=LB
.param LB3=LB

.param L1=Phi0/(4*IC*Ic0)
.param L2=(Phi0/(2*B1*Ic0))/2
.param L3=L2
.param L4=Phi0/(4*IC*Ic0)
.param L5=L3
.param L6=L4

.param LP1=LP
.param LP2=LP
.param LP3=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 8 9 jjmit  area=B3 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 10 pwl(0 0 5p IB3)

LB1 3 1 1.712E-012 
LB2 7 5 2.279E-012 
LB3 10 8 2.858E-012 

L1 a 1 2.062E-012 
L2 1 4 2.06E-012 
L3 5 4 2.079E-012 
L4 5 q0 2.081E-012 
L5 4 8 2.076E-012 
L6 8 q1 2.086E-012 

LP1 2 0 4.263E-013 
LP2 6 0 3.75E-013 
LP3 9 0 4.312E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 8 108 RB3  
LRB3 108 0 LRB3 

.ends
