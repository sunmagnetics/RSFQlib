* Author: L. Schindler
* Version: 2.1
* Last modification date: 28 April 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

*$Ports 			a clk q
.subckt LSmitll_NOTT a clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param RD=1.36
.param LB=0.2p
.param Lptl=2p
.param LP=0.5p

.param B1=1.26
.param B2=1.42
.param B3=1.72 
.param B4=1.22
.param B5=0.77
.param B6=1.40
.param B7=2.5
.param B8=2
.param B9=1.35
.param B10=1.04 
.param B11=1.41
.param B12=2.5

.param IB1=173u
.param IB2=123u
.param IB3=230u
.param IB4=112u
.param IB5=112u
.param IB6=108u
.param IB7=187u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB

.param L1=Lptl
.param L2=4.4718p
.param L3=2.6117p
.param L4=1.1676p
.param L5=2.6532p 
.param L7=3.1681p
.param L8=0.86946p
.param L9=Lptl
.param L10=2.5468p
.param L11=2.1566p
.param L12=0.99180p
.param L13=3.286p
.param L14=6.5962p
.param L15=0.42413p
.param L16=2.2847p
.param L17=0.49986p 
.param L18=0.28417p
.param L19=7.3651p
.param L20=0.74611p
.param L21=4.5195p
.param L22=Lptl

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12

.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet

B1 2 3 jjmit area=B1
B2 6 7 jjmit area=B2
B3 10 12 jjmit area=B3
B4 15 14 jjmit area=B4
B5 15 31 jjmit area=B5
B6 17 18 jjmit area=B6
B7 21 22 jjmit area=B7
B8 25 26 jjmit area=B8
B9 29 30 jjmit area=B9
B10 32 33 jjmit area=B10
B11 36 37 jjmit area=B11
B12 38 40 jjmit area=B12

IB1 0 5 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
IB3 0 20 pwl(0 0 5p IB3)
IB4 0 24 pwl(0 0 5p IB4)
IB5 0 28 pwl(0 0 5p IB5)
IB6 0 35 pwl(0 0 5p IB6)
IB7 0 39 pwl(0 0 5p IB7)

L1 a 2 L1
L2 2 4 L2
L3 4 6 L3
L4 6 8 L4
L5 8 10 L5
L7 10 13 L7
L8 10 14 L8
L9 clk 17 L9
L10 17 19 L10 
L11 19 21 L11
L12 21 23 L12
L13 23 25 L13
L14 25 27 L14
L15 27 15 L15
L16 25 29 L16
L17 30 31 L17
L18 30 32 L18
L19 32 34 L19
L20 34 36 L20
L21 36 38 L21
L22 38 41 L22

RN 13 0 3.54
RD 41 q RD

LB1 4 5 LB1
LB2 8 9 LB2
LB3 19 20 LB3
LB4 23 24 LB4
LB5 27 28 LB5
LB6 34 35 LB6
LB7 38 39 LB7

LP1 3 0 LP
LP2 7 0 LP
LP3 12 0 LP
LP6 18 0 LP
LP7 22 0 LP
LP8 26 0 LP
LP10 33 0 LP
LP11 37 0 LP
LP12 40 0 LP

RB1 2 102 RB1
LRB1 102 0 LRB1
RB2 6 106 RB2
LRB2 106 0 LRB2
RB3 10 110 RB3
LRB3 110 0 LRB3
RB4 14 114 RB4
LRB4 114 15 LRB4
RB5 15 115 RB5
LRB5 115 31 LRB5
RB6 17 117 RB6
LRB6 117 0 LRB6
RB7 21 121 RB7
LRB7 121 0 LRB7
RB8 25 125 RB8
LRB8 125 0 LRB8
RB9 29 129 RB9
LRB9 129 30 LRB9
RB10 32 132 RB10
LRB10 132 0 LRB10
RB11 36 136 RB11
LRB11 136 0 LRB11
RB12 38 138 RB12
LRB12 138 0 LRB12
.ends