* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/18.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 16 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Tessa Hall, 19775539@sun.ac.za

*$ports 	a	b	clk	q
.subckt THmitll_OR2T a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param ICreceive=1.6
.param ICtrans=2.5
.param LB=2p
.param BiasCoef=0.7
.param Lptl=2p
.param RD=1.36

.param B1=1.6
.param B2=1.28
.param B3=1.65
.param B4=1.25
.param B5=1.6
.param B6=1.28
.param B7=1.65
.param B8=1.25
.param B9=1.67
.param B10=1.95
.param B11=1.6
.param B12=1.59
.param B13=1.44
.param B14=2.09
.param B15=2.5

.param IB1=112u
.param IB2=156u
.param IB3=112u
.param IB4=156u
.param IB5=210u
.param IB6=176u
.param IB7=242u
.param IB8=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param LB8=LB

.param L1=Lptl
.param L2=6.7019p
.param L3=6.2519p
.param L4=0.7723p
.param L5=Lptl
.param L6=6.7019p
.param L7=6.2519p
.param L8=0.7723p
.param L9=4.6089p
.param L10=7.7141p
.param L11=Lptl
.param L12=2.7407p
.param L13=3.4070p
.param L14=4.5212p
.param L15=4.5560p
.param L16=Lptl

.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LP5=LP
.param LP6=LP
.param LP7=LP
.param LP10=LP
.param LP11=LP
.param LP12=LP
.param LP14=LP
.param LP15=LP

.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11   
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet+LP 
.param LRB6=(RB6/Rsheet)*Lsheet+LP
.param LRB7=(RB7/Rsheet)*Lsheet+LP 
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet+LP
.param LRB12=(RB12/Rsheet)*Lsheet+LP
.param LRB13=(RB13/Rsheet)*Lsheet
.param LRB14=(RB14/Rsheet)*Lsheet+LP
.param LRB15=(RB15/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
B4 7 9 jjmit  area=B4 
B5 11 12 jjmit  area=B5 
B6 14 15 jjmit  area=B6 
B7 17 18 jjmit  area=B7 
B8 17 19 jjmit  area=B8 
B9 21 22 jjmit  area=B9 
B10 22 23 jjmit  area=B10 
B11 26 27 jjmit  area=B11 
B12 30 31 jjmit  area=B12 
B13 32 25 jjmit  area=B13 
B14 25 33 jjmit  area=B14 
B15 34 35 jjmit  area=B15 

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 6 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 16 pwl(0 0 5p IB4)
IB5 0 20 pwl(0 0 5p IB5)
IB6 0 24 pwl(0 0 5p IB6)
IB7 0 29 pwl(0 0 5p IB7)
IB8 0 36 pwl(0 0 5p IB8)

LB1 3 1 4.448E-012 
LB2 6 4 2.203E-012 
LB3 13 11 4.442E-012 
LB4 16 14 2.187E-012 
LB5 20 10 3.603E-012 
LB6 24 22 1.443E-012 
LB7 29 28 1.069E-012 
LB8 36 34 8.669E-013 

L1 a 1 1.444E-012 
L2 1 4 6.665E-012 
L3 4 7 6.254E-012 
L4 9 10 7.702E-013 
L5 b 11 1.443E-012 
L6 11 14 6.656E-012 
L7 14 17 6.244E-012 
L8 19 10 7.773E-013 
L9 10 21 4.573E-012 
L10 22 25 7.702E-012 
L11 clk 26 1.282E-012 
L12 26 28 2.735E-012 
L13 28 30 3.418E-012 
L14 30 32 4.48E-012 
L15 25 34 4.553E-012 
L16 34 37 8.104E-013 

RD 37 q RD  

LP1 2 0 4.195E-013 
LP2 5 0 5.813E-013 
LP3 8 0 4.455E-013 
LP5 12 0 4.193E-013 
LP6 15 0 5.831E-013 
LP7 18 0 4.774E-013 
LP10 23 0 4.819E-013 
LP11 27 0 3.541E-013 
LP12 31 0 4.657E-013 
LP14 33 0 4.19E-013 
LP15 35 0 3.333E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3 
RB4 7 109 RB4  
LRB4 109 9 LRB4 
RB5 11 111 RB5  
LRB5 111 0 LRB5 
RB6 14 114 RB6  
LRB6 114 0 LRB6 
RB7 17 117 RB7  
LRB7 117 0 LRB7 
RB8 17 119 RB8  
LRB8 119 19 LRB8 
RB9 21 121 RB9  
LRB9 121 22 LRB9 
RB10 22 122 RB10  
LRB10 122 0 LRB10 
RB11 26 126 RB11  
LRB11 126 0 LRB11 
RB12 30 130 RB12  
LRB12 130 0 LRB12 
RB13 32 132 RB13  
LRB13 132 25 LRB13 
RB14 25 125 RB14  
LRB14 125 0 LRB14 
RB15 34 134 RB15  
LRB15 134 0 LRB15 

.ends
