* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

*$Ports 			a q
.subckt LSmitll_PTLRX_SFQDC a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
B00 103 108 jjmit area=1
B01 104 110 jjmit area=1
B02 105 112 jjmit area=1
I00 0 106 pwl(0 0 5p 155u)
L00 106 107 0.2p
L01 a 103 0.2p
L02 103 107 4.3p
L03 107 104 4.6p
L04 104 105 5p
L05 105 5001 2.3p
L06 108 0 0.34p
L07 109 0 0.5p
L08 110 0 0.06p
L09 111 0 1p
L010 112 0 0.03p
L011 113 0 1p
R00 103 109 6.859904418
R01 104 111 6.859904418
R02 105 113 6.859904418

.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param B1=3.25
.param B2=2.00
.param B3=1.50
.param B4=3.00
.param B5=1.75
.param B6=1.50
.param B7=1.50
.param B8=2.00
.param L1=1.522p
.param L3=0.827p
.param L4=1.12884p
.param L5=1.11098p
.param L6=5.940p
.param L7=3.216p
.param L10=0.215p
.param L13=3.699p
.param L17=1.510p
.param L18=2.010p
.param L19=0.954p
.param L4b=0.178p
.param LB1=(RB1/Rsheet)*Lsheet
.param LB2=(RB2/Rsheet)*Lsheet
.param LB3=(RB3/Rsheet)*Lsheet
.param LB4=(RB4/Rsheet)*Lsheet
.param LB5=(RB5/Rsheet)*Lsheet
.param LB6=(RB6/Rsheet)*Lsheet
.param LB7=(RB7/Rsheet)*Lsheet
.param LB8=(RB8/Rsheet)*Lsheet
.param LP1=0.140p
.param LP4=0.524p
.param LP5=0.516p
.param LP7=0.086p
.param LP8=0.226p
.param LR1=0.91p
.param R1=0.375
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param IB1=280u
.param IB2=150u
.param IB3=220u
.param IB4=80u
B1 8 20 jjmit area=B1
B2 12 13 jjmit area=B2
B3 3 4 jjmit area=B3
B4 13 29 jjmit area=B4
B5 5 16 jjmit area=B5
B6 6 7 jjmit area=B6
B7 10 22 jjmit area=B7
B8 11 24 jjmit area=B8
IB1 0 8 pwl(0 0 5p IB1)
IB2 0 4 pwl(0 0 5p IB2)
IB3 0 7 pwl(0 0 5p IB3)
IB4 0 18 pwl(0 0 5p IB4)
L1 5001 8 L1
L3 8 17 L3
L4 3 17 L4
L5 17 12 L5
L6 5 9 L6
L7 9 13 L7
L10 9 6 L10
L13 10 18 L13
L17 11 q L17
L18 18 11 L18
L19 7 10 L19
L4b 4 5 L4b
LB1 8 21 LB1
LB2 12 27 LB2
LB3 3 14 LB3
LB4 13 28 LB4
LB5 5 15 LB5
LB6 6 19 LB6
LB7 10 23 LB7
LB8 11 25 LB8
LP1 20 0 LP1
LP4 29 0 LP4
LP5 16 0 LP5
LP7 22 0 LP7
LP8 24 0 LP8
LR1 9 26 LR1
R1 26 0 R1
RB1 21 0 RB1
RB2 27 13 RB2
RB3 14 4 RB3
RB4 28 0 RB4
RB5 15 0 RB5
RB6 19 7 RB6
RB7 23 0 RB7
RB8 25 0 RB8
.ends