* Author: L. Schindler
* Version: 2.1
* Last modification date: 3 June 2021
* Last modification by: L. Schindler

* Copyright (c) 2018-2021 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, lschindler@sun.ac.za

* The cell is not designed to be connected directly to passive transmission lines

*$Ports		a		clk		q
.subckt LSmitll_DFF	  a	clk q	
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.70

.param B1=IC
.param B2=IC/1.4
.param B3=IC
.param B4=IC
.param B5=IC/1.4
.param B6=IC
.param B7=IC

.param IB1=BiasCoef*Ic0*B1         
.param IB2=Ic0*Ic          
.param IB3=BiasCoef*Ic0*B6             
.param IB4=BiasCoef*Ic0*B7         

.param L1=Phi0/(4*IC*Ic0)               
.param L2=Phi0/(2*B1*Ic0)         
.param L3=Phi0/(B3*Ic0)       
.param L4=Phi0/(2*B6*Ic0)      
.param L5=Phi0/(4*IC*Ic0)     
.param L6=Phi0/(2*B4*Ic0)       
.param L7=Phi0/(4*B7*Ic0)         
.param LB1=LB           
.param LB2=LB          
.param LB3=LB           
.param LB4=LB         
.param LP1=LP         
.param LP3=LP          
.param LP4=LP         
.param LP6=LP          
.param LP7=LP          
.param RB1=B0Rs/B1       
.param RB2=B0Rs/B2       
.param RB3=B0Rs/B3          
.param RB4=B0Rs/B4         
.param RB5=B0Rs/B5         
.param RB6=B0Rs/B6          
.param RB7=B0Rs/B7
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet
.param LRB4=(RB4/Rsheet)*Lsheet
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet

B1 1 2 jjmit area=B1
B2 4 5 jjmit area=B2
B3 5 6 jjmit area=B3
B4 8 9 jjmit area=B4
B5 10 8 jjmit area=B5
B6 11 12 jjmit area=B6
B7 14 15 jjmit area=B7

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 13 pwl(0 0 5p IB3)
IB4 0 16 pwl(0 0 5p IB4)

LB1 3 1 LB1
LB2 7 5 LB2
LB3 11 13 LB3
LB4 16 14 LB4

L1 a 1 L1
L2 1 4 L2
L3 5 8 L3
L4 10 11 L4
L5 clk 11 L5
L6 8 14 L6
L7 14 q L7

LP1 2 0 LP1    
LP3 6 0 LP3    
LP4 9 0 LP4    
LP6 12 0 LP6    
LP7 15 0 LP7    

RB1 1 101 RB1
LRB1 101 0 LRB1
RB2 4 104 RB2
LRB2 104 5 LRB2
RB3 5 105 RB3
LRB3 105 0 LRB3
RB4 8 108 RB4
LRB4 108 0 LRB4
RB5 10 110 RB5
LRB5 110 8 LRB5
RB6 11 111 RB6
LRB6 111 0 LRB6
RB7 14 114 RB7
LRB7 114 0 LRB7
.ends