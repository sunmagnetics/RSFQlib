* Back-annotated simulation file written by InductEx v.6.1.52 on 2022/08/09.
* Author: L. Schindler
* Version: 3.0
* Last modification date: 4 August 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

* The cell is not designed to be connected directly to passive transmission lines.

*$Ports 	a	b	clk	q
.subckt THmitll_AND2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7

.param B1=2.5
.param B2=1.60
.param B3=1.94
.param B4=1.57
.param B5=1.25
.param B6=1.25
.param B7=2.5
.param B8=1.60
.param B9=1.94
.param B10=1.57
.param B11=1.25
.param B12=1.25
.param B13=2.5
.param B14=1.71
.param B15=2.5

.param IB1=175u
.param IB2=162u
.param IB3=175u
.param IB4=162u
.param IB5=175u
.param IB6=124u
.param IB7=175u

.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB

.param L1=1.8843p
.param L2=4.2266p
.param L3=9.6820p
.param L4=0.9913p
.param L5=2.5745p
.param L6=1.8843p
.param L7=4.2266p
.param L8=9.6820p
.param L9=0.9913p
.param L10=2.5745p
.param L11=1.5293p
.param L12=2.6230p
.param L13=0.7965p
.param L14=0.7671p
.param L15=1.2144p

.param LP1=LP
.param LP3=LP
.param LP4=LP
.param LP7=LP
.param LP9=LP
.param LP10=LP
.param LP13=LP
.param LP14=LP
.param LP15=LP

.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15

.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet+LP
.param LRB14=(RB14/Rsheet)*Lsheet+LP
.param LRB15=(RB15/Rsheet)*Lsheet+LP

B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 5 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 8 10 jjmit  area=B5 
B6 12 13 jjmit  area=B6 
B7 14 15 jjmit  area=B7 
B8 17 18 jjmit  area=B8 
B9 18 19 jjmit  area=B9 
B10 21 22 jjmit  area=B10 
B11 21 23 jjmit  area=B11 
B12 24 13 jjmit  area=B12 
B13 25 26 jjmit  area=B13 
B14 28 29 jjmit  area=B14 
B15 31 32 jjmit  area=B15

IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 27 pwl(0 0 5p IB5)
IB6 0 30 pwl(0 0 5p IB6)
IB7 0 33 pwl(0 0 5p IB7)

LB1 3 1 1.032E-012 
LB2 7 5 3.135E-012 
LB3 16 14 1.016E-012 
LB4 20 18 3.19E-012 
LB5 27 25 1.708E-012 
LB6 30 28 6.363E-013 
LB7 33 31 7.55E-013 

L1 a 1 1.874E-012 
L2 1 4 4.249E-012 
L3 5 8 9.672E-012 
L4 10 11 9.976E-013 
L5 8 12 2.561E-012 
L6 b 14 1.875E-012 
L7 14 17 4.233E-012 
L8 18 21 9.691E-012 
L9 11 23 9.928E-013 
L10 21 24 2.556E-012 
L11 clk 25 1.531E-012 
L12 25 28 2.626E-012 
L13 28 11 7.973E-013 
L14 13 31 7.691E-013 
L15 31 q 1.217E-012 

LP1 2 0 3.464E-013 
LP3 6 0 6.827E-013 
LP4 0 9 4.723E-013 
LP7 15 0 3.484E-013 
LP9 19 0 6.81E-013 
LP10 22 0 4.756E-013 
LP13 26 0 3.392E-013 
LP14 29 0 3.972E-013 
LP15 32 0 3.699E-013 

RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 5 LRB2 
RB3 5 105 RB3  
LRB3 105 0 LRB3 
RB4 108 8 RB4  
LRB4 0 108 LRB4 
RB5 8 110 RB5  
LRB5 110 10 LRB5 
RB6 12 112 RB6  
LRB6 112 13 LRB6 
RB7 14 114 RB7  
LRB7 114 0 LRB7 
RB8 17 117 RB8  
LRB8 117 18 LRB8 
RB9 18 118 RB9  
LRB9 118 0 LRB9 
RB10 21 121 RB10  
LRB10 121 0 LRB10 
RB11 123 21 RB11  
LRB11 23 123 LRB11 
RB12 24 124 RB12  
LRB12 124 13 LRB12 
RB13 25 125 RB13  
LRB13 125 0 LRB13 
RB14 28 128 RB14  
LRB14 128 0 LRB14 
RB15 31 131 RB15  
LRB15 131 0 LRB15 

.ends
