* Manually Generated Testbench
* Author: T. Hall
* Version: 3.0
* Last modification date: 22 July 2022
* Last modification by: T. Hall

* Copyright (c) 2018-2022 Lieze Schindler, Tessa Hall, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

* For questions about the library, contact Tessa Hall, 19775539@sun.ac.za.

*-----------------------
* SINK CELL: RESISTOR
*-----------------------

.subckt sinkcell out
rsink out 0 2
.ends

*-----------------------
*  LOAD OUT CELL: JTL
*-----------------------

.subckt THmitll_JTL a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7
.param B1=IC
.param B2=IC
.param IB1=(B1+B2)*Ic0*BiasCoef
.param LB1=LB
.param L1=Phi0/(4*B1*Ic0)
.param L2=Phi0/(4*B1*Ic0)
.param L3=Phi0/(4*B2*Ic0)
.param L4=Phi0/(4*B2*Ic0)
.param LP1=LP
.param LP2=LP
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
B1 1 2 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
IB1 0 4 pwl(0 0 5p IB1)
LB1 4 3 2.336E-012 
L1 a 1 2.07E-012 
L2 1 3 2.088E-012 
L3 3 5 2.082E-012 
L4 5 q 2.072E-012 
LP1 2 0 3.137E-013 
LP2 6 0 3.123E-013 
RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
.ends

*-----------------------
*  TEST DEVICE: DCSFQ
*-----------------------

.subckt THmitll_DCSFQ a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7
.param B1=2.25
.param B2=2.25
.param B3=IC
.param IB1=275u
.param IB2=B3*Ic0*BiasCoef
.param LB1=LB
.param LB2=LB
.param L1=1p
.param L2=3.9p
.param L3=0.6p
.param L4=1.1p
.param L5=4.5p
.param L6=Phi0/(4*IC*Ic0)
.param LP2=LP
.param LP3=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
B1 2 3 jjmit  area=B1 
B2 5 6 jjmit  area=B2 
B3 7 8 jjmit  area=B3 
IB1 0 4 pwl(0 0 5p IB1)
IB2 0 9 pwl(0 0 5p IB2)
LB1 4 3 2.825E-012 
LB2 9 7 2.942E-012 
L1 a 1 1.672E-012 
L2 1 0 3.901E-012 
L3 1 2 5.953E-013 
L4 3 5 1.1E-012 
L5 5 7 4.542E-012 
L6 7 q 2.012E-012 
LP2 6 0 3.924E-013 
LP3 8 0 3.841E-013 
RB1 2 102 RB1  
LRB1 102 3 LRB1 
RB2 5 105 RB2  
LRB2 105 0 LRB2 
RB3 7 107 RB3  
LRB3 107 0 LRB3
.ends

*-----------------------
*        CONTROL
*-----------------------

I_a 0 a pulse(0 600u 20p 2p 2p 1p 100p)
XDUT THmitll_DCSFQ a q
XLOADOUT THmitll_JTL q out
XRout  sinkcell	out

.tran 0.025p 1000p 0
.print i(L1.XDUT) i(L6.XDUT) p(B3.XDUT) p(B1.XLOADOUT)
.end