* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 3.0
* Last modification date: 23 August 2022
* Last modification by: T. Hall

.control
	back-annotate THmitll_ALWAYS0_SYNC_v3p0_base.cir
.endc

L1 a 1 2.0678p [L1]
L2 1 4 4.1357p [L2]
L3 clk 5 2.0678p [L3]
L4 5 8 4.1357p [L4]
L5 9 10 4.1357p [L5]
L6 10 q 2.0678p [L6]

LB1 1 3 [LB1]
LB2 5 7 [LB2]
LB3 10 12 [LB3]

LP1 2 0 [LP1]
LP2 6 0 [LP2]
LP3 11 0 [LP3]

* Ports
P1 a 0
P2 clk 0
P3 q 0

J1 1 2 250u
J2 5 6 250u
J3 10 11 250u

PB1 3 0
PB2 7 0
PB3 12 0

PR1 4 0
PR2 8 0
PR3 9 0
.end